library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity fft_pt2048 is
    GENERIC (
        ctrl_start     : INTEGER := 0
    );
    PORT (
        tmp_first_stage_re_out, tmp_first_stage_im_out: OUT STD_LOGIC_VECTOR(2047 DOWNTO 0);
        tmp_mul_re_out, tmp_mul_im_out : OUT STD_LOGIC_VECTOR(2047 DOWNTO 0);

        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        bypass         : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        ctrl           : IN STD_LOGIC;

        data_re_in     : IN STD_LOGIC_VECTOR(2047 DOWNTO 0);
        data_im_in     : IN STD_LOGIC_VECTOR(2047 DOWNTO 0);

        data_re_out    : OUT STD_LOGIC_VECTOR(2047 DOWNTO 0);
        data_im_out    : OUT STD_LOGIC_VECTOR(2047 DOWNTO 0)
    );
end fft_pt2048;

architecture Behavioral of fft_pt2048 is

component fft_pt32 is
    GENERIC (
        ctrl_start     : INTEGER
    );
    PORT (
        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        bypass         : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        ctrl_delay     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

        data_re_in     : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        data_im_in     : IN STD_LOGIC_VECTOR(31 DOWNTO 0);

        data_re_out    : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        data_im_out    : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
end component;

component fft_pt64 is
    GENERIC (
        ctrl_start       : INTEGER
    );
    PORT (
        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        bypass         : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
        ctrl_delay     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

        data_re_in     : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
        data_im_in     : IN STD_LOGIC_VECTOR(63 DOWNTO 0);

        data_re_out     : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
        data_im_out     : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
    );
end component;

component complex_multiplier is
    GENERIC (
        ctrl_start       : INTEGER
    );
    PORT (
        clk              : IN STD_LOGIC;
        rst              : IN STD_LOGIC;
        ce               : IN STD_LOGIC;
        bypass           : IN STD_LOGIC;
        ctrl_delay       : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_in       : IN STD_LOGIC;
        data_im_in       : IN STD_LOGIC;
        re_multiplicator : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        im_multiplicator : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_out      : OUT STD_LOGIC;
        data_im_out      : OUT STD_LOGIC
    );
end component;

component multiplier_mul1 IS
    GENERIC (
        ctrl_start : INTEGER := 0
    );
    PORT (
        clk             : IN STD_LOGIC;
        rst             : IN STD_LOGIC;
        ce              : IN STD_LOGIC;
        bypass          : IN STD_LOGIC;
        ctrl_delay      : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_in      : IN STD_LOGIC;
        data_im_in      : IN STD_LOGIC;
        data_re_out     : OUT STD_LOGIC;
        data_im_out     : OUT STD_LOGIC
    );
END component;

component multiplier_mulminusj IS
    GENERIC (
        ctrl_start : INTEGER := 0
    );
    PORT (
        clk             : IN STD_LOGIC;
        rst             : IN STD_LOGIC;
        ce              : IN STD_LOGIC;
        bypass          : IN STD_LOGIC;
        ctrl_delay      : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_in      : IN STD_LOGIC;
        data_im_in      : IN STD_LOGIC;
        data_re_out     : OUT STD_LOGIC;
        data_im_out     : OUT STD_LOGIC
    );
END component;

COMPONENT Dff_regN_Nout IS
    GENERIC (N : INTEGER);
    PORT (  
        D      : IN STD_LOGIC;
        clk    : IN STD_LOGIC;
        Q      : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        QN     : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0)
    );
END COMPONENT;

signal first_stage_re_out, first_stage_im_out: STD_LOGIC_VECTOR(2047 DOWNTO 0);
signal mul_re_out, mul_im_out : STD_LOGIC_VECTOR(2047 DOWNTO 0);

SIGNAL ctrl_delay : STD_LOGIC_VECTOR(15 DOWNTO 0);

begin
    --- create ctrl_delay signal IN top module
    ctrl_delay(0) <= ctrl;
    --- buffer for ctrl
    UDFF_CTRL : Dff_regN_Nout
    GENERIC MAP(
        N => 15
    )
    PORT MAP(
        D           => ctrl, 
        clk         => clk, 
        Q           => ctrl_delay(15 DOWNTO 1)
    );


    tmp_first_stage_re_out <= first_stage_re_out;
    tmp_first_stage_im_out <= first_stage_im_out;
    tmp_mul_re_out <= mul_re_out;
    tmp_mul_im_out <= mul_im_out;

    --- left-hand-side processors
    ULFFT_PT32_0 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(0),
            data_re_in(1) => data_re_in(64),
            data_re_in(2) => data_re_in(128),
            data_re_in(3) => data_re_in(192),
            data_re_in(4) => data_re_in(256),
            data_re_in(5) => data_re_in(320),
            data_re_in(6) => data_re_in(384),
            data_re_in(7) => data_re_in(448),
            data_re_in(8) => data_re_in(512),
            data_re_in(9) => data_re_in(576),
            data_re_in(10) => data_re_in(640),
            data_re_in(11) => data_re_in(704),
            data_re_in(12) => data_re_in(768),
            data_re_in(13) => data_re_in(832),
            data_re_in(14) => data_re_in(896),
            data_re_in(15) => data_re_in(960),
            data_re_in(16) => data_re_in(1024),
            data_re_in(17) => data_re_in(1088),
            data_re_in(18) => data_re_in(1152),
            data_re_in(19) => data_re_in(1216),
            data_re_in(20) => data_re_in(1280),
            data_re_in(21) => data_re_in(1344),
            data_re_in(22) => data_re_in(1408),
            data_re_in(23) => data_re_in(1472),
            data_re_in(24) => data_re_in(1536),
            data_re_in(25) => data_re_in(1600),
            data_re_in(26) => data_re_in(1664),
            data_re_in(27) => data_re_in(1728),
            data_re_in(28) => data_re_in(1792),
            data_re_in(29) => data_re_in(1856),
            data_re_in(30) => data_re_in(1920),
            data_re_in(31) => data_re_in(1984),
            data_im_in(0) => data_im_in(0),
            data_im_in(1) => data_im_in(64),
            data_im_in(2) => data_im_in(128),
            data_im_in(3) => data_im_in(192),
            data_im_in(4) => data_im_in(256),
            data_im_in(5) => data_im_in(320),
            data_im_in(6) => data_im_in(384),
            data_im_in(7) => data_im_in(448),
            data_im_in(8) => data_im_in(512),
            data_im_in(9) => data_im_in(576),
            data_im_in(10) => data_im_in(640),
            data_im_in(11) => data_im_in(704),
            data_im_in(12) => data_im_in(768),
            data_im_in(13) => data_im_in(832),
            data_im_in(14) => data_im_in(896),
            data_im_in(15) => data_im_in(960),
            data_im_in(16) => data_im_in(1024),
            data_im_in(17) => data_im_in(1088),
            data_im_in(18) => data_im_in(1152),
            data_im_in(19) => data_im_in(1216),
            data_im_in(20) => data_im_in(1280),
            data_im_in(21) => data_im_in(1344),
            data_im_in(22) => data_im_in(1408),
            data_im_in(23) => data_im_in(1472),
            data_im_in(24) => data_im_in(1536),
            data_im_in(25) => data_im_in(1600),
            data_im_in(26) => data_im_in(1664),
            data_im_in(27) => data_im_in(1728),
            data_im_in(28) => data_im_in(1792),
            data_im_in(29) => data_im_in(1856),
            data_im_in(30) => data_im_in(1920),
            data_im_in(31) => data_im_in(1984),
            data_re_out(0) => first_stage_re_out(0),
            data_re_out(1) => first_stage_re_out(64),
            data_re_out(2) => first_stage_re_out(128),
            data_re_out(3) => first_stage_re_out(192),
            data_re_out(4) => first_stage_re_out(256),
            data_re_out(5) => first_stage_re_out(320),
            data_re_out(6) => first_stage_re_out(384),
            data_re_out(7) => first_stage_re_out(448),
            data_re_out(8) => first_stage_re_out(512),
            data_re_out(9) => first_stage_re_out(576),
            data_re_out(10) => first_stage_re_out(640),
            data_re_out(11) => first_stage_re_out(704),
            data_re_out(12) => first_stage_re_out(768),
            data_re_out(13) => first_stage_re_out(832),
            data_re_out(14) => first_stage_re_out(896),
            data_re_out(15) => first_stage_re_out(960),
            data_re_out(16) => first_stage_re_out(1024),
            data_re_out(17) => first_stage_re_out(1088),
            data_re_out(18) => first_stage_re_out(1152),
            data_re_out(19) => first_stage_re_out(1216),
            data_re_out(20) => first_stage_re_out(1280),
            data_re_out(21) => first_stage_re_out(1344),
            data_re_out(22) => first_stage_re_out(1408),
            data_re_out(23) => first_stage_re_out(1472),
            data_re_out(24) => first_stage_re_out(1536),
            data_re_out(25) => first_stage_re_out(1600),
            data_re_out(26) => first_stage_re_out(1664),
            data_re_out(27) => first_stage_re_out(1728),
            data_re_out(28) => first_stage_re_out(1792),
            data_re_out(29) => first_stage_re_out(1856),
            data_re_out(30) => first_stage_re_out(1920),
            data_re_out(31) => first_stage_re_out(1984),
            data_im_out(0) => first_stage_im_out(0),
            data_im_out(1) => first_stage_im_out(64),
            data_im_out(2) => first_stage_im_out(128),
            data_im_out(3) => first_stage_im_out(192),
            data_im_out(4) => first_stage_im_out(256),
            data_im_out(5) => first_stage_im_out(320),
            data_im_out(6) => first_stage_im_out(384),
            data_im_out(7) => first_stage_im_out(448),
            data_im_out(8) => first_stage_im_out(512),
            data_im_out(9) => first_stage_im_out(576),
            data_im_out(10) => first_stage_im_out(640),
            data_im_out(11) => first_stage_im_out(704),
            data_im_out(12) => first_stage_im_out(768),
            data_im_out(13) => first_stage_im_out(832),
            data_im_out(14) => first_stage_im_out(896),
            data_im_out(15) => first_stage_im_out(960),
            data_im_out(16) => first_stage_im_out(1024),
            data_im_out(17) => first_stage_im_out(1088),
            data_im_out(18) => first_stage_im_out(1152),
            data_im_out(19) => first_stage_im_out(1216),
            data_im_out(20) => first_stage_im_out(1280),
            data_im_out(21) => first_stage_im_out(1344),
            data_im_out(22) => first_stage_im_out(1408),
            data_im_out(23) => first_stage_im_out(1472),
            data_im_out(24) => first_stage_im_out(1536),
            data_im_out(25) => first_stage_im_out(1600),
            data_im_out(26) => first_stage_im_out(1664),
            data_im_out(27) => first_stage_im_out(1728),
            data_im_out(28) => first_stage_im_out(1792),
            data_im_out(29) => first_stage_im_out(1856),
            data_im_out(30) => first_stage_im_out(1920),
            data_im_out(31) => first_stage_im_out(1984)
        );

    ULFFT_PT32_1 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(1),
            data_re_in(1) => data_re_in(65),
            data_re_in(2) => data_re_in(129),
            data_re_in(3) => data_re_in(193),
            data_re_in(4) => data_re_in(257),
            data_re_in(5) => data_re_in(321),
            data_re_in(6) => data_re_in(385),
            data_re_in(7) => data_re_in(449),
            data_re_in(8) => data_re_in(513),
            data_re_in(9) => data_re_in(577),
            data_re_in(10) => data_re_in(641),
            data_re_in(11) => data_re_in(705),
            data_re_in(12) => data_re_in(769),
            data_re_in(13) => data_re_in(833),
            data_re_in(14) => data_re_in(897),
            data_re_in(15) => data_re_in(961),
            data_re_in(16) => data_re_in(1025),
            data_re_in(17) => data_re_in(1089),
            data_re_in(18) => data_re_in(1153),
            data_re_in(19) => data_re_in(1217),
            data_re_in(20) => data_re_in(1281),
            data_re_in(21) => data_re_in(1345),
            data_re_in(22) => data_re_in(1409),
            data_re_in(23) => data_re_in(1473),
            data_re_in(24) => data_re_in(1537),
            data_re_in(25) => data_re_in(1601),
            data_re_in(26) => data_re_in(1665),
            data_re_in(27) => data_re_in(1729),
            data_re_in(28) => data_re_in(1793),
            data_re_in(29) => data_re_in(1857),
            data_re_in(30) => data_re_in(1921),
            data_re_in(31) => data_re_in(1985),
            data_im_in(0) => data_im_in(1),
            data_im_in(1) => data_im_in(65),
            data_im_in(2) => data_im_in(129),
            data_im_in(3) => data_im_in(193),
            data_im_in(4) => data_im_in(257),
            data_im_in(5) => data_im_in(321),
            data_im_in(6) => data_im_in(385),
            data_im_in(7) => data_im_in(449),
            data_im_in(8) => data_im_in(513),
            data_im_in(9) => data_im_in(577),
            data_im_in(10) => data_im_in(641),
            data_im_in(11) => data_im_in(705),
            data_im_in(12) => data_im_in(769),
            data_im_in(13) => data_im_in(833),
            data_im_in(14) => data_im_in(897),
            data_im_in(15) => data_im_in(961),
            data_im_in(16) => data_im_in(1025),
            data_im_in(17) => data_im_in(1089),
            data_im_in(18) => data_im_in(1153),
            data_im_in(19) => data_im_in(1217),
            data_im_in(20) => data_im_in(1281),
            data_im_in(21) => data_im_in(1345),
            data_im_in(22) => data_im_in(1409),
            data_im_in(23) => data_im_in(1473),
            data_im_in(24) => data_im_in(1537),
            data_im_in(25) => data_im_in(1601),
            data_im_in(26) => data_im_in(1665),
            data_im_in(27) => data_im_in(1729),
            data_im_in(28) => data_im_in(1793),
            data_im_in(29) => data_im_in(1857),
            data_im_in(30) => data_im_in(1921),
            data_im_in(31) => data_im_in(1985),
            data_re_out(0) => first_stage_re_out(1),
            data_re_out(1) => first_stage_re_out(65),
            data_re_out(2) => first_stage_re_out(129),
            data_re_out(3) => first_stage_re_out(193),
            data_re_out(4) => first_stage_re_out(257),
            data_re_out(5) => first_stage_re_out(321),
            data_re_out(6) => first_stage_re_out(385),
            data_re_out(7) => first_stage_re_out(449),
            data_re_out(8) => first_stage_re_out(513),
            data_re_out(9) => first_stage_re_out(577),
            data_re_out(10) => first_stage_re_out(641),
            data_re_out(11) => first_stage_re_out(705),
            data_re_out(12) => first_stage_re_out(769),
            data_re_out(13) => first_stage_re_out(833),
            data_re_out(14) => first_stage_re_out(897),
            data_re_out(15) => first_stage_re_out(961),
            data_re_out(16) => first_stage_re_out(1025),
            data_re_out(17) => first_stage_re_out(1089),
            data_re_out(18) => first_stage_re_out(1153),
            data_re_out(19) => first_stage_re_out(1217),
            data_re_out(20) => first_stage_re_out(1281),
            data_re_out(21) => first_stage_re_out(1345),
            data_re_out(22) => first_stage_re_out(1409),
            data_re_out(23) => first_stage_re_out(1473),
            data_re_out(24) => first_stage_re_out(1537),
            data_re_out(25) => first_stage_re_out(1601),
            data_re_out(26) => first_stage_re_out(1665),
            data_re_out(27) => first_stage_re_out(1729),
            data_re_out(28) => first_stage_re_out(1793),
            data_re_out(29) => first_stage_re_out(1857),
            data_re_out(30) => first_stage_re_out(1921),
            data_re_out(31) => first_stage_re_out(1985),
            data_im_out(0) => first_stage_im_out(1),
            data_im_out(1) => first_stage_im_out(65),
            data_im_out(2) => first_stage_im_out(129),
            data_im_out(3) => first_stage_im_out(193),
            data_im_out(4) => first_stage_im_out(257),
            data_im_out(5) => first_stage_im_out(321),
            data_im_out(6) => first_stage_im_out(385),
            data_im_out(7) => first_stage_im_out(449),
            data_im_out(8) => first_stage_im_out(513),
            data_im_out(9) => first_stage_im_out(577),
            data_im_out(10) => first_stage_im_out(641),
            data_im_out(11) => first_stage_im_out(705),
            data_im_out(12) => first_stage_im_out(769),
            data_im_out(13) => first_stage_im_out(833),
            data_im_out(14) => first_stage_im_out(897),
            data_im_out(15) => first_stage_im_out(961),
            data_im_out(16) => first_stage_im_out(1025),
            data_im_out(17) => first_stage_im_out(1089),
            data_im_out(18) => first_stage_im_out(1153),
            data_im_out(19) => first_stage_im_out(1217),
            data_im_out(20) => first_stage_im_out(1281),
            data_im_out(21) => first_stage_im_out(1345),
            data_im_out(22) => first_stage_im_out(1409),
            data_im_out(23) => first_stage_im_out(1473),
            data_im_out(24) => first_stage_im_out(1537),
            data_im_out(25) => first_stage_im_out(1601),
            data_im_out(26) => first_stage_im_out(1665),
            data_im_out(27) => first_stage_im_out(1729),
            data_im_out(28) => first_stage_im_out(1793),
            data_im_out(29) => first_stage_im_out(1857),
            data_im_out(30) => first_stage_im_out(1921),
            data_im_out(31) => first_stage_im_out(1985)
        );

    ULFFT_PT32_2 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(2),
            data_re_in(1) => data_re_in(66),
            data_re_in(2) => data_re_in(130),
            data_re_in(3) => data_re_in(194),
            data_re_in(4) => data_re_in(258),
            data_re_in(5) => data_re_in(322),
            data_re_in(6) => data_re_in(386),
            data_re_in(7) => data_re_in(450),
            data_re_in(8) => data_re_in(514),
            data_re_in(9) => data_re_in(578),
            data_re_in(10) => data_re_in(642),
            data_re_in(11) => data_re_in(706),
            data_re_in(12) => data_re_in(770),
            data_re_in(13) => data_re_in(834),
            data_re_in(14) => data_re_in(898),
            data_re_in(15) => data_re_in(962),
            data_re_in(16) => data_re_in(1026),
            data_re_in(17) => data_re_in(1090),
            data_re_in(18) => data_re_in(1154),
            data_re_in(19) => data_re_in(1218),
            data_re_in(20) => data_re_in(1282),
            data_re_in(21) => data_re_in(1346),
            data_re_in(22) => data_re_in(1410),
            data_re_in(23) => data_re_in(1474),
            data_re_in(24) => data_re_in(1538),
            data_re_in(25) => data_re_in(1602),
            data_re_in(26) => data_re_in(1666),
            data_re_in(27) => data_re_in(1730),
            data_re_in(28) => data_re_in(1794),
            data_re_in(29) => data_re_in(1858),
            data_re_in(30) => data_re_in(1922),
            data_re_in(31) => data_re_in(1986),
            data_im_in(0) => data_im_in(2),
            data_im_in(1) => data_im_in(66),
            data_im_in(2) => data_im_in(130),
            data_im_in(3) => data_im_in(194),
            data_im_in(4) => data_im_in(258),
            data_im_in(5) => data_im_in(322),
            data_im_in(6) => data_im_in(386),
            data_im_in(7) => data_im_in(450),
            data_im_in(8) => data_im_in(514),
            data_im_in(9) => data_im_in(578),
            data_im_in(10) => data_im_in(642),
            data_im_in(11) => data_im_in(706),
            data_im_in(12) => data_im_in(770),
            data_im_in(13) => data_im_in(834),
            data_im_in(14) => data_im_in(898),
            data_im_in(15) => data_im_in(962),
            data_im_in(16) => data_im_in(1026),
            data_im_in(17) => data_im_in(1090),
            data_im_in(18) => data_im_in(1154),
            data_im_in(19) => data_im_in(1218),
            data_im_in(20) => data_im_in(1282),
            data_im_in(21) => data_im_in(1346),
            data_im_in(22) => data_im_in(1410),
            data_im_in(23) => data_im_in(1474),
            data_im_in(24) => data_im_in(1538),
            data_im_in(25) => data_im_in(1602),
            data_im_in(26) => data_im_in(1666),
            data_im_in(27) => data_im_in(1730),
            data_im_in(28) => data_im_in(1794),
            data_im_in(29) => data_im_in(1858),
            data_im_in(30) => data_im_in(1922),
            data_im_in(31) => data_im_in(1986),
            data_re_out(0) => first_stage_re_out(2),
            data_re_out(1) => first_stage_re_out(66),
            data_re_out(2) => first_stage_re_out(130),
            data_re_out(3) => first_stage_re_out(194),
            data_re_out(4) => first_stage_re_out(258),
            data_re_out(5) => first_stage_re_out(322),
            data_re_out(6) => first_stage_re_out(386),
            data_re_out(7) => first_stage_re_out(450),
            data_re_out(8) => first_stage_re_out(514),
            data_re_out(9) => first_stage_re_out(578),
            data_re_out(10) => first_stage_re_out(642),
            data_re_out(11) => first_stage_re_out(706),
            data_re_out(12) => first_stage_re_out(770),
            data_re_out(13) => first_stage_re_out(834),
            data_re_out(14) => first_stage_re_out(898),
            data_re_out(15) => first_stage_re_out(962),
            data_re_out(16) => first_stage_re_out(1026),
            data_re_out(17) => first_stage_re_out(1090),
            data_re_out(18) => first_stage_re_out(1154),
            data_re_out(19) => first_stage_re_out(1218),
            data_re_out(20) => first_stage_re_out(1282),
            data_re_out(21) => first_stage_re_out(1346),
            data_re_out(22) => first_stage_re_out(1410),
            data_re_out(23) => first_stage_re_out(1474),
            data_re_out(24) => first_stage_re_out(1538),
            data_re_out(25) => first_stage_re_out(1602),
            data_re_out(26) => first_stage_re_out(1666),
            data_re_out(27) => first_stage_re_out(1730),
            data_re_out(28) => first_stage_re_out(1794),
            data_re_out(29) => first_stage_re_out(1858),
            data_re_out(30) => first_stage_re_out(1922),
            data_re_out(31) => first_stage_re_out(1986),
            data_im_out(0) => first_stage_im_out(2),
            data_im_out(1) => first_stage_im_out(66),
            data_im_out(2) => first_stage_im_out(130),
            data_im_out(3) => first_stage_im_out(194),
            data_im_out(4) => first_stage_im_out(258),
            data_im_out(5) => first_stage_im_out(322),
            data_im_out(6) => first_stage_im_out(386),
            data_im_out(7) => first_stage_im_out(450),
            data_im_out(8) => first_stage_im_out(514),
            data_im_out(9) => first_stage_im_out(578),
            data_im_out(10) => first_stage_im_out(642),
            data_im_out(11) => first_stage_im_out(706),
            data_im_out(12) => first_stage_im_out(770),
            data_im_out(13) => first_stage_im_out(834),
            data_im_out(14) => first_stage_im_out(898),
            data_im_out(15) => first_stage_im_out(962),
            data_im_out(16) => first_stage_im_out(1026),
            data_im_out(17) => first_stage_im_out(1090),
            data_im_out(18) => first_stage_im_out(1154),
            data_im_out(19) => first_stage_im_out(1218),
            data_im_out(20) => first_stage_im_out(1282),
            data_im_out(21) => first_stage_im_out(1346),
            data_im_out(22) => first_stage_im_out(1410),
            data_im_out(23) => first_stage_im_out(1474),
            data_im_out(24) => first_stage_im_out(1538),
            data_im_out(25) => first_stage_im_out(1602),
            data_im_out(26) => first_stage_im_out(1666),
            data_im_out(27) => first_stage_im_out(1730),
            data_im_out(28) => first_stage_im_out(1794),
            data_im_out(29) => first_stage_im_out(1858),
            data_im_out(30) => first_stage_im_out(1922),
            data_im_out(31) => first_stage_im_out(1986)
        );

    ULFFT_PT32_3 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(3),
            data_re_in(1) => data_re_in(67),
            data_re_in(2) => data_re_in(131),
            data_re_in(3) => data_re_in(195),
            data_re_in(4) => data_re_in(259),
            data_re_in(5) => data_re_in(323),
            data_re_in(6) => data_re_in(387),
            data_re_in(7) => data_re_in(451),
            data_re_in(8) => data_re_in(515),
            data_re_in(9) => data_re_in(579),
            data_re_in(10) => data_re_in(643),
            data_re_in(11) => data_re_in(707),
            data_re_in(12) => data_re_in(771),
            data_re_in(13) => data_re_in(835),
            data_re_in(14) => data_re_in(899),
            data_re_in(15) => data_re_in(963),
            data_re_in(16) => data_re_in(1027),
            data_re_in(17) => data_re_in(1091),
            data_re_in(18) => data_re_in(1155),
            data_re_in(19) => data_re_in(1219),
            data_re_in(20) => data_re_in(1283),
            data_re_in(21) => data_re_in(1347),
            data_re_in(22) => data_re_in(1411),
            data_re_in(23) => data_re_in(1475),
            data_re_in(24) => data_re_in(1539),
            data_re_in(25) => data_re_in(1603),
            data_re_in(26) => data_re_in(1667),
            data_re_in(27) => data_re_in(1731),
            data_re_in(28) => data_re_in(1795),
            data_re_in(29) => data_re_in(1859),
            data_re_in(30) => data_re_in(1923),
            data_re_in(31) => data_re_in(1987),
            data_im_in(0) => data_im_in(3),
            data_im_in(1) => data_im_in(67),
            data_im_in(2) => data_im_in(131),
            data_im_in(3) => data_im_in(195),
            data_im_in(4) => data_im_in(259),
            data_im_in(5) => data_im_in(323),
            data_im_in(6) => data_im_in(387),
            data_im_in(7) => data_im_in(451),
            data_im_in(8) => data_im_in(515),
            data_im_in(9) => data_im_in(579),
            data_im_in(10) => data_im_in(643),
            data_im_in(11) => data_im_in(707),
            data_im_in(12) => data_im_in(771),
            data_im_in(13) => data_im_in(835),
            data_im_in(14) => data_im_in(899),
            data_im_in(15) => data_im_in(963),
            data_im_in(16) => data_im_in(1027),
            data_im_in(17) => data_im_in(1091),
            data_im_in(18) => data_im_in(1155),
            data_im_in(19) => data_im_in(1219),
            data_im_in(20) => data_im_in(1283),
            data_im_in(21) => data_im_in(1347),
            data_im_in(22) => data_im_in(1411),
            data_im_in(23) => data_im_in(1475),
            data_im_in(24) => data_im_in(1539),
            data_im_in(25) => data_im_in(1603),
            data_im_in(26) => data_im_in(1667),
            data_im_in(27) => data_im_in(1731),
            data_im_in(28) => data_im_in(1795),
            data_im_in(29) => data_im_in(1859),
            data_im_in(30) => data_im_in(1923),
            data_im_in(31) => data_im_in(1987),
            data_re_out(0) => first_stage_re_out(3),
            data_re_out(1) => first_stage_re_out(67),
            data_re_out(2) => first_stage_re_out(131),
            data_re_out(3) => first_stage_re_out(195),
            data_re_out(4) => first_stage_re_out(259),
            data_re_out(5) => first_stage_re_out(323),
            data_re_out(6) => first_stage_re_out(387),
            data_re_out(7) => first_stage_re_out(451),
            data_re_out(8) => first_stage_re_out(515),
            data_re_out(9) => first_stage_re_out(579),
            data_re_out(10) => first_stage_re_out(643),
            data_re_out(11) => first_stage_re_out(707),
            data_re_out(12) => first_stage_re_out(771),
            data_re_out(13) => first_stage_re_out(835),
            data_re_out(14) => first_stage_re_out(899),
            data_re_out(15) => first_stage_re_out(963),
            data_re_out(16) => first_stage_re_out(1027),
            data_re_out(17) => first_stage_re_out(1091),
            data_re_out(18) => first_stage_re_out(1155),
            data_re_out(19) => first_stage_re_out(1219),
            data_re_out(20) => first_stage_re_out(1283),
            data_re_out(21) => first_stage_re_out(1347),
            data_re_out(22) => first_stage_re_out(1411),
            data_re_out(23) => first_stage_re_out(1475),
            data_re_out(24) => first_stage_re_out(1539),
            data_re_out(25) => first_stage_re_out(1603),
            data_re_out(26) => first_stage_re_out(1667),
            data_re_out(27) => first_stage_re_out(1731),
            data_re_out(28) => first_stage_re_out(1795),
            data_re_out(29) => first_stage_re_out(1859),
            data_re_out(30) => first_stage_re_out(1923),
            data_re_out(31) => first_stage_re_out(1987),
            data_im_out(0) => first_stage_im_out(3),
            data_im_out(1) => first_stage_im_out(67),
            data_im_out(2) => first_stage_im_out(131),
            data_im_out(3) => first_stage_im_out(195),
            data_im_out(4) => first_stage_im_out(259),
            data_im_out(5) => first_stage_im_out(323),
            data_im_out(6) => first_stage_im_out(387),
            data_im_out(7) => first_stage_im_out(451),
            data_im_out(8) => first_stage_im_out(515),
            data_im_out(9) => first_stage_im_out(579),
            data_im_out(10) => first_stage_im_out(643),
            data_im_out(11) => first_stage_im_out(707),
            data_im_out(12) => first_stage_im_out(771),
            data_im_out(13) => first_stage_im_out(835),
            data_im_out(14) => first_stage_im_out(899),
            data_im_out(15) => first_stage_im_out(963),
            data_im_out(16) => first_stage_im_out(1027),
            data_im_out(17) => first_stage_im_out(1091),
            data_im_out(18) => first_stage_im_out(1155),
            data_im_out(19) => first_stage_im_out(1219),
            data_im_out(20) => first_stage_im_out(1283),
            data_im_out(21) => first_stage_im_out(1347),
            data_im_out(22) => first_stage_im_out(1411),
            data_im_out(23) => first_stage_im_out(1475),
            data_im_out(24) => first_stage_im_out(1539),
            data_im_out(25) => first_stage_im_out(1603),
            data_im_out(26) => first_stage_im_out(1667),
            data_im_out(27) => first_stage_im_out(1731),
            data_im_out(28) => first_stage_im_out(1795),
            data_im_out(29) => first_stage_im_out(1859),
            data_im_out(30) => first_stage_im_out(1923),
            data_im_out(31) => first_stage_im_out(1987)
        );

    ULFFT_PT32_4 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(4),
            data_re_in(1) => data_re_in(68),
            data_re_in(2) => data_re_in(132),
            data_re_in(3) => data_re_in(196),
            data_re_in(4) => data_re_in(260),
            data_re_in(5) => data_re_in(324),
            data_re_in(6) => data_re_in(388),
            data_re_in(7) => data_re_in(452),
            data_re_in(8) => data_re_in(516),
            data_re_in(9) => data_re_in(580),
            data_re_in(10) => data_re_in(644),
            data_re_in(11) => data_re_in(708),
            data_re_in(12) => data_re_in(772),
            data_re_in(13) => data_re_in(836),
            data_re_in(14) => data_re_in(900),
            data_re_in(15) => data_re_in(964),
            data_re_in(16) => data_re_in(1028),
            data_re_in(17) => data_re_in(1092),
            data_re_in(18) => data_re_in(1156),
            data_re_in(19) => data_re_in(1220),
            data_re_in(20) => data_re_in(1284),
            data_re_in(21) => data_re_in(1348),
            data_re_in(22) => data_re_in(1412),
            data_re_in(23) => data_re_in(1476),
            data_re_in(24) => data_re_in(1540),
            data_re_in(25) => data_re_in(1604),
            data_re_in(26) => data_re_in(1668),
            data_re_in(27) => data_re_in(1732),
            data_re_in(28) => data_re_in(1796),
            data_re_in(29) => data_re_in(1860),
            data_re_in(30) => data_re_in(1924),
            data_re_in(31) => data_re_in(1988),
            data_im_in(0) => data_im_in(4),
            data_im_in(1) => data_im_in(68),
            data_im_in(2) => data_im_in(132),
            data_im_in(3) => data_im_in(196),
            data_im_in(4) => data_im_in(260),
            data_im_in(5) => data_im_in(324),
            data_im_in(6) => data_im_in(388),
            data_im_in(7) => data_im_in(452),
            data_im_in(8) => data_im_in(516),
            data_im_in(9) => data_im_in(580),
            data_im_in(10) => data_im_in(644),
            data_im_in(11) => data_im_in(708),
            data_im_in(12) => data_im_in(772),
            data_im_in(13) => data_im_in(836),
            data_im_in(14) => data_im_in(900),
            data_im_in(15) => data_im_in(964),
            data_im_in(16) => data_im_in(1028),
            data_im_in(17) => data_im_in(1092),
            data_im_in(18) => data_im_in(1156),
            data_im_in(19) => data_im_in(1220),
            data_im_in(20) => data_im_in(1284),
            data_im_in(21) => data_im_in(1348),
            data_im_in(22) => data_im_in(1412),
            data_im_in(23) => data_im_in(1476),
            data_im_in(24) => data_im_in(1540),
            data_im_in(25) => data_im_in(1604),
            data_im_in(26) => data_im_in(1668),
            data_im_in(27) => data_im_in(1732),
            data_im_in(28) => data_im_in(1796),
            data_im_in(29) => data_im_in(1860),
            data_im_in(30) => data_im_in(1924),
            data_im_in(31) => data_im_in(1988),
            data_re_out(0) => first_stage_re_out(4),
            data_re_out(1) => first_stage_re_out(68),
            data_re_out(2) => first_stage_re_out(132),
            data_re_out(3) => first_stage_re_out(196),
            data_re_out(4) => first_stage_re_out(260),
            data_re_out(5) => first_stage_re_out(324),
            data_re_out(6) => first_stage_re_out(388),
            data_re_out(7) => first_stage_re_out(452),
            data_re_out(8) => first_stage_re_out(516),
            data_re_out(9) => first_stage_re_out(580),
            data_re_out(10) => first_stage_re_out(644),
            data_re_out(11) => first_stage_re_out(708),
            data_re_out(12) => first_stage_re_out(772),
            data_re_out(13) => first_stage_re_out(836),
            data_re_out(14) => first_stage_re_out(900),
            data_re_out(15) => first_stage_re_out(964),
            data_re_out(16) => first_stage_re_out(1028),
            data_re_out(17) => first_stage_re_out(1092),
            data_re_out(18) => first_stage_re_out(1156),
            data_re_out(19) => first_stage_re_out(1220),
            data_re_out(20) => first_stage_re_out(1284),
            data_re_out(21) => first_stage_re_out(1348),
            data_re_out(22) => first_stage_re_out(1412),
            data_re_out(23) => first_stage_re_out(1476),
            data_re_out(24) => first_stage_re_out(1540),
            data_re_out(25) => first_stage_re_out(1604),
            data_re_out(26) => first_stage_re_out(1668),
            data_re_out(27) => first_stage_re_out(1732),
            data_re_out(28) => first_stage_re_out(1796),
            data_re_out(29) => first_stage_re_out(1860),
            data_re_out(30) => first_stage_re_out(1924),
            data_re_out(31) => first_stage_re_out(1988),
            data_im_out(0) => first_stage_im_out(4),
            data_im_out(1) => first_stage_im_out(68),
            data_im_out(2) => first_stage_im_out(132),
            data_im_out(3) => first_stage_im_out(196),
            data_im_out(4) => first_stage_im_out(260),
            data_im_out(5) => first_stage_im_out(324),
            data_im_out(6) => first_stage_im_out(388),
            data_im_out(7) => first_stage_im_out(452),
            data_im_out(8) => first_stage_im_out(516),
            data_im_out(9) => first_stage_im_out(580),
            data_im_out(10) => first_stage_im_out(644),
            data_im_out(11) => first_stage_im_out(708),
            data_im_out(12) => first_stage_im_out(772),
            data_im_out(13) => first_stage_im_out(836),
            data_im_out(14) => first_stage_im_out(900),
            data_im_out(15) => first_stage_im_out(964),
            data_im_out(16) => first_stage_im_out(1028),
            data_im_out(17) => first_stage_im_out(1092),
            data_im_out(18) => first_stage_im_out(1156),
            data_im_out(19) => first_stage_im_out(1220),
            data_im_out(20) => first_stage_im_out(1284),
            data_im_out(21) => first_stage_im_out(1348),
            data_im_out(22) => first_stage_im_out(1412),
            data_im_out(23) => first_stage_im_out(1476),
            data_im_out(24) => first_stage_im_out(1540),
            data_im_out(25) => first_stage_im_out(1604),
            data_im_out(26) => first_stage_im_out(1668),
            data_im_out(27) => first_stage_im_out(1732),
            data_im_out(28) => first_stage_im_out(1796),
            data_im_out(29) => first_stage_im_out(1860),
            data_im_out(30) => first_stage_im_out(1924),
            data_im_out(31) => first_stage_im_out(1988)
        );

    ULFFT_PT32_5 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(5),
            data_re_in(1) => data_re_in(69),
            data_re_in(2) => data_re_in(133),
            data_re_in(3) => data_re_in(197),
            data_re_in(4) => data_re_in(261),
            data_re_in(5) => data_re_in(325),
            data_re_in(6) => data_re_in(389),
            data_re_in(7) => data_re_in(453),
            data_re_in(8) => data_re_in(517),
            data_re_in(9) => data_re_in(581),
            data_re_in(10) => data_re_in(645),
            data_re_in(11) => data_re_in(709),
            data_re_in(12) => data_re_in(773),
            data_re_in(13) => data_re_in(837),
            data_re_in(14) => data_re_in(901),
            data_re_in(15) => data_re_in(965),
            data_re_in(16) => data_re_in(1029),
            data_re_in(17) => data_re_in(1093),
            data_re_in(18) => data_re_in(1157),
            data_re_in(19) => data_re_in(1221),
            data_re_in(20) => data_re_in(1285),
            data_re_in(21) => data_re_in(1349),
            data_re_in(22) => data_re_in(1413),
            data_re_in(23) => data_re_in(1477),
            data_re_in(24) => data_re_in(1541),
            data_re_in(25) => data_re_in(1605),
            data_re_in(26) => data_re_in(1669),
            data_re_in(27) => data_re_in(1733),
            data_re_in(28) => data_re_in(1797),
            data_re_in(29) => data_re_in(1861),
            data_re_in(30) => data_re_in(1925),
            data_re_in(31) => data_re_in(1989),
            data_im_in(0) => data_im_in(5),
            data_im_in(1) => data_im_in(69),
            data_im_in(2) => data_im_in(133),
            data_im_in(3) => data_im_in(197),
            data_im_in(4) => data_im_in(261),
            data_im_in(5) => data_im_in(325),
            data_im_in(6) => data_im_in(389),
            data_im_in(7) => data_im_in(453),
            data_im_in(8) => data_im_in(517),
            data_im_in(9) => data_im_in(581),
            data_im_in(10) => data_im_in(645),
            data_im_in(11) => data_im_in(709),
            data_im_in(12) => data_im_in(773),
            data_im_in(13) => data_im_in(837),
            data_im_in(14) => data_im_in(901),
            data_im_in(15) => data_im_in(965),
            data_im_in(16) => data_im_in(1029),
            data_im_in(17) => data_im_in(1093),
            data_im_in(18) => data_im_in(1157),
            data_im_in(19) => data_im_in(1221),
            data_im_in(20) => data_im_in(1285),
            data_im_in(21) => data_im_in(1349),
            data_im_in(22) => data_im_in(1413),
            data_im_in(23) => data_im_in(1477),
            data_im_in(24) => data_im_in(1541),
            data_im_in(25) => data_im_in(1605),
            data_im_in(26) => data_im_in(1669),
            data_im_in(27) => data_im_in(1733),
            data_im_in(28) => data_im_in(1797),
            data_im_in(29) => data_im_in(1861),
            data_im_in(30) => data_im_in(1925),
            data_im_in(31) => data_im_in(1989),
            data_re_out(0) => first_stage_re_out(5),
            data_re_out(1) => first_stage_re_out(69),
            data_re_out(2) => first_stage_re_out(133),
            data_re_out(3) => first_stage_re_out(197),
            data_re_out(4) => first_stage_re_out(261),
            data_re_out(5) => first_stage_re_out(325),
            data_re_out(6) => first_stage_re_out(389),
            data_re_out(7) => first_stage_re_out(453),
            data_re_out(8) => first_stage_re_out(517),
            data_re_out(9) => first_stage_re_out(581),
            data_re_out(10) => first_stage_re_out(645),
            data_re_out(11) => first_stage_re_out(709),
            data_re_out(12) => first_stage_re_out(773),
            data_re_out(13) => first_stage_re_out(837),
            data_re_out(14) => first_stage_re_out(901),
            data_re_out(15) => first_stage_re_out(965),
            data_re_out(16) => first_stage_re_out(1029),
            data_re_out(17) => first_stage_re_out(1093),
            data_re_out(18) => first_stage_re_out(1157),
            data_re_out(19) => first_stage_re_out(1221),
            data_re_out(20) => first_stage_re_out(1285),
            data_re_out(21) => first_stage_re_out(1349),
            data_re_out(22) => first_stage_re_out(1413),
            data_re_out(23) => first_stage_re_out(1477),
            data_re_out(24) => first_stage_re_out(1541),
            data_re_out(25) => first_stage_re_out(1605),
            data_re_out(26) => first_stage_re_out(1669),
            data_re_out(27) => first_stage_re_out(1733),
            data_re_out(28) => first_stage_re_out(1797),
            data_re_out(29) => first_stage_re_out(1861),
            data_re_out(30) => first_stage_re_out(1925),
            data_re_out(31) => first_stage_re_out(1989),
            data_im_out(0) => first_stage_im_out(5),
            data_im_out(1) => first_stage_im_out(69),
            data_im_out(2) => first_stage_im_out(133),
            data_im_out(3) => first_stage_im_out(197),
            data_im_out(4) => first_stage_im_out(261),
            data_im_out(5) => first_stage_im_out(325),
            data_im_out(6) => first_stage_im_out(389),
            data_im_out(7) => first_stage_im_out(453),
            data_im_out(8) => first_stage_im_out(517),
            data_im_out(9) => first_stage_im_out(581),
            data_im_out(10) => first_stage_im_out(645),
            data_im_out(11) => first_stage_im_out(709),
            data_im_out(12) => first_stage_im_out(773),
            data_im_out(13) => first_stage_im_out(837),
            data_im_out(14) => first_stage_im_out(901),
            data_im_out(15) => first_stage_im_out(965),
            data_im_out(16) => first_stage_im_out(1029),
            data_im_out(17) => first_stage_im_out(1093),
            data_im_out(18) => first_stage_im_out(1157),
            data_im_out(19) => first_stage_im_out(1221),
            data_im_out(20) => first_stage_im_out(1285),
            data_im_out(21) => first_stage_im_out(1349),
            data_im_out(22) => first_stage_im_out(1413),
            data_im_out(23) => first_stage_im_out(1477),
            data_im_out(24) => first_stage_im_out(1541),
            data_im_out(25) => first_stage_im_out(1605),
            data_im_out(26) => first_stage_im_out(1669),
            data_im_out(27) => first_stage_im_out(1733),
            data_im_out(28) => first_stage_im_out(1797),
            data_im_out(29) => first_stage_im_out(1861),
            data_im_out(30) => first_stage_im_out(1925),
            data_im_out(31) => first_stage_im_out(1989)
        );

    ULFFT_PT32_6 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(6),
            data_re_in(1) => data_re_in(70),
            data_re_in(2) => data_re_in(134),
            data_re_in(3) => data_re_in(198),
            data_re_in(4) => data_re_in(262),
            data_re_in(5) => data_re_in(326),
            data_re_in(6) => data_re_in(390),
            data_re_in(7) => data_re_in(454),
            data_re_in(8) => data_re_in(518),
            data_re_in(9) => data_re_in(582),
            data_re_in(10) => data_re_in(646),
            data_re_in(11) => data_re_in(710),
            data_re_in(12) => data_re_in(774),
            data_re_in(13) => data_re_in(838),
            data_re_in(14) => data_re_in(902),
            data_re_in(15) => data_re_in(966),
            data_re_in(16) => data_re_in(1030),
            data_re_in(17) => data_re_in(1094),
            data_re_in(18) => data_re_in(1158),
            data_re_in(19) => data_re_in(1222),
            data_re_in(20) => data_re_in(1286),
            data_re_in(21) => data_re_in(1350),
            data_re_in(22) => data_re_in(1414),
            data_re_in(23) => data_re_in(1478),
            data_re_in(24) => data_re_in(1542),
            data_re_in(25) => data_re_in(1606),
            data_re_in(26) => data_re_in(1670),
            data_re_in(27) => data_re_in(1734),
            data_re_in(28) => data_re_in(1798),
            data_re_in(29) => data_re_in(1862),
            data_re_in(30) => data_re_in(1926),
            data_re_in(31) => data_re_in(1990),
            data_im_in(0) => data_im_in(6),
            data_im_in(1) => data_im_in(70),
            data_im_in(2) => data_im_in(134),
            data_im_in(3) => data_im_in(198),
            data_im_in(4) => data_im_in(262),
            data_im_in(5) => data_im_in(326),
            data_im_in(6) => data_im_in(390),
            data_im_in(7) => data_im_in(454),
            data_im_in(8) => data_im_in(518),
            data_im_in(9) => data_im_in(582),
            data_im_in(10) => data_im_in(646),
            data_im_in(11) => data_im_in(710),
            data_im_in(12) => data_im_in(774),
            data_im_in(13) => data_im_in(838),
            data_im_in(14) => data_im_in(902),
            data_im_in(15) => data_im_in(966),
            data_im_in(16) => data_im_in(1030),
            data_im_in(17) => data_im_in(1094),
            data_im_in(18) => data_im_in(1158),
            data_im_in(19) => data_im_in(1222),
            data_im_in(20) => data_im_in(1286),
            data_im_in(21) => data_im_in(1350),
            data_im_in(22) => data_im_in(1414),
            data_im_in(23) => data_im_in(1478),
            data_im_in(24) => data_im_in(1542),
            data_im_in(25) => data_im_in(1606),
            data_im_in(26) => data_im_in(1670),
            data_im_in(27) => data_im_in(1734),
            data_im_in(28) => data_im_in(1798),
            data_im_in(29) => data_im_in(1862),
            data_im_in(30) => data_im_in(1926),
            data_im_in(31) => data_im_in(1990),
            data_re_out(0) => first_stage_re_out(6),
            data_re_out(1) => first_stage_re_out(70),
            data_re_out(2) => first_stage_re_out(134),
            data_re_out(3) => first_stage_re_out(198),
            data_re_out(4) => first_stage_re_out(262),
            data_re_out(5) => first_stage_re_out(326),
            data_re_out(6) => first_stage_re_out(390),
            data_re_out(7) => first_stage_re_out(454),
            data_re_out(8) => first_stage_re_out(518),
            data_re_out(9) => first_stage_re_out(582),
            data_re_out(10) => first_stage_re_out(646),
            data_re_out(11) => first_stage_re_out(710),
            data_re_out(12) => first_stage_re_out(774),
            data_re_out(13) => first_stage_re_out(838),
            data_re_out(14) => first_stage_re_out(902),
            data_re_out(15) => first_stage_re_out(966),
            data_re_out(16) => first_stage_re_out(1030),
            data_re_out(17) => first_stage_re_out(1094),
            data_re_out(18) => first_stage_re_out(1158),
            data_re_out(19) => first_stage_re_out(1222),
            data_re_out(20) => first_stage_re_out(1286),
            data_re_out(21) => first_stage_re_out(1350),
            data_re_out(22) => first_stage_re_out(1414),
            data_re_out(23) => first_stage_re_out(1478),
            data_re_out(24) => first_stage_re_out(1542),
            data_re_out(25) => first_stage_re_out(1606),
            data_re_out(26) => first_stage_re_out(1670),
            data_re_out(27) => first_stage_re_out(1734),
            data_re_out(28) => first_stage_re_out(1798),
            data_re_out(29) => first_stage_re_out(1862),
            data_re_out(30) => first_stage_re_out(1926),
            data_re_out(31) => first_stage_re_out(1990),
            data_im_out(0) => first_stage_im_out(6),
            data_im_out(1) => first_stage_im_out(70),
            data_im_out(2) => first_stage_im_out(134),
            data_im_out(3) => first_stage_im_out(198),
            data_im_out(4) => first_stage_im_out(262),
            data_im_out(5) => first_stage_im_out(326),
            data_im_out(6) => first_stage_im_out(390),
            data_im_out(7) => first_stage_im_out(454),
            data_im_out(8) => first_stage_im_out(518),
            data_im_out(9) => first_stage_im_out(582),
            data_im_out(10) => first_stage_im_out(646),
            data_im_out(11) => first_stage_im_out(710),
            data_im_out(12) => first_stage_im_out(774),
            data_im_out(13) => first_stage_im_out(838),
            data_im_out(14) => first_stage_im_out(902),
            data_im_out(15) => first_stage_im_out(966),
            data_im_out(16) => first_stage_im_out(1030),
            data_im_out(17) => first_stage_im_out(1094),
            data_im_out(18) => first_stage_im_out(1158),
            data_im_out(19) => first_stage_im_out(1222),
            data_im_out(20) => first_stage_im_out(1286),
            data_im_out(21) => first_stage_im_out(1350),
            data_im_out(22) => first_stage_im_out(1414),
            data_im_out(23) => first_stage_im_out(1478),
            data_im_out(24) => first_stage_im_out(1542),
            data_im_out(25) => first_stage_im_out(1606),
            data_im_out(26) => first_stage_im_out(1670),
            data_im_out(27) => first_stage_im_out(1734),
            data_im_out(28) => first_stage_im_out(1798),
            data_im_out(29) => first_stage_im_out(1862),
            data_im_out(30) => first_stage_im_out(1926),
            data_im_out(31) => first_stage_im_out(1990)
        );

    ULFFT_PT32_7 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(7),
            data_re_in(1) => data_re_in(71),
            data_re_in(2) => data_re_in(135),
            data_re_in(3) => data_re_in(199),
            data_re_in(4) => data_re_in(263),
            data_re_in(5) => data_re_in(327),
            data_re_in(6) => data_re_in(391),
            data_re_in(7) => data_re_in(455),
            data_re_in(8) => data_re_in(519),
            data_re_in(9) => data_re_in(583),
            data_re_in(10) => data_re_in(647),
            data_re_in(11) => data_re_in(711),
            data_re_in(12) => data_re_in(775),
            data_re_in(13) => data_re_in(839),
            data_re_in(14) => data_re_in(903),
            data_re_in(15) => data_re_in(967),
            data_re_in(16) => data_re_in(1031),
            data_re_in(17) => data_re_in(1095),
            data_re_in(18) => data_re_in(1159),
            data_re_in(19) => data_re_in(1223),
            data_re_in(20) => data_re_in(1287),
            data_re_in(21) => data_re_in(1351),
            data_re_in(22) => data_re_in(1415),
            data_re_in(23) => data_re_in(1479),
            data_re_in(24) => data_re_in(1543),
            data_re_in(25) => data_re_in(1607),
            data_re_in(26) => data_re_in(1671),
            data_re_in(27) => data_re_in(1735),
            data_re_in(28) => data_re_in(1799),
            data_re_in(29) => data_re_in(1863),
            data_re_in(30) => data_re_in(1927),
            data_re_in(31) => data_re_in(1991),
            data_im_in(0) => data_im_in(7),
            data_im_in(1) => data_im_in(71),
            data_im_in(2) => data_im_in(135),
            data_im_in(3) => data_im_in(199),
            data_im_in(4) => data_im_in(263),
            data_im_in(5) => data_im_in(327),
            data_im_in(6) => data_im_in(391),
            data_im_in(7) => data_im_in(455),
            data_im_in(8) => data_im_in(519),
            data_im_in(9) => data_im_in(583),
            data_im_in(10) => data_im_in(647),
            data_im_in(11) => data_im_in(711),
            data_im_in(12) => data_im_in(775),
            data_im_in(13) => data_im_in(839),
            data_im_in(14) => data_im_in(903),
            data_im_in(15) => data_im_in(967),
            data_im_in(16) => data_im_in(1031),
            data_im_in(17) => data_im_in(1095),
            data_im_in(18) => data_im_in(1159),
            data_im_in(19) => data_im_in(1223),
            data_im_in(20) => data_im_in(1287),
            data_im_in(21) => data_im_in(1351),
            data_im_in(22) => data_im_in(1415),
            data_im_in(23) => data_im_in(1479),
            data_im_in(24) => data_im_in(1543),
            data_im_in(25) => data_im_in(1607),
            data_im_in(26) => data_im_in(1671),
            data_im_in(27) => data_im_in(1735),
            data_im_in(28) => data_im_in(1799),
            data_im_in(29) => data_im_in(1863),
            data_im_in(30) => data_im_in(1927),
            data_im_in(31) => data_im_in(1991),
            data_re_out(0) => first_stage_re_out(7),
            data_re_out(1) => first_stage_re_out(71),
            data_re_out(2) => first_stage_re_out(135),
            data_re_out(3) => first_stage_re_out(199),
            data_re_out(4) => first_stage_re_out(263),
            data_re_out(5) => first_stage_re_out(327),
            data_re_out(6) => first_stage_re_out(391),
            data_re_out(7) => first_stage_re_out(455),
            data_re_out(8) => first_stage_re_out(519),
            data_re_out(9) => first_stage_re_out(583),
            data_re_out(10) => first_stage_re_out(647),
            data_re_out(11) => first_stage_re_out(711),
            data_re_out(12) => first_stage_re_out(775),
            data_re_out(13) => first_stage_re_out(839),
            data_re_out(14) => first_stage_re_out(903),
            data_re_out(15) => first_stage_re_out(967),
            data_re_out(16) => first_stage_re_out(1031),
            data_re_out(17) => first_stage_re_out(1095),
            data_re_out(18) => first_stage_re_out(1159),
            data_re_out(19) => first_stage_re_out(1223),
            data_re_out(20) => first_stage_re_out(1287),
            data_re_out(21) => first_stage_re_out(1351),
            data_re_out(22) => first_stage_re_out(1415),
            data_re_out(23) => first_stage_re_out(1479),
            data_re_out(24) => first_stage_re_out(1543),
            data_re_out(25) => first_stage_re_out(1607),
            data_re_out(26) => first_stage_re_out(1671),
            data_re_out(27) => first_stage_re_out(1735),
            data_re_out(28) => first_stage_re_out(1799),
            data_re_out(29) => first_stage_re_out(1863),
            data_re_out(30) => first_stage_re_out(1927),
            data_re_out(31) => first_stage_re_out(1991),
            data_im_out(0) => first_stage_im_out(7),
            data_im_out(1) => first_stage_im_out(71),
            data_im_out(2) => first_stage_im_out(135),
            data_im_out(3) => first_stage_im_out(199),
            data_im_out(4) => first_stage_im_out(263),
            data_im_out(5) => first_stage_im_out(327),
            data_im_out(6) => first_stage_im_out(391),
            data_im_out(7) => first_stage_im_out(455),
            data_im_out(8) => first_stage_im_out(519),
            data_im_out(9) => first_stage_im_out(583),
            data_im_out(10) => first_stage_im_out(647),
            data_im_out(11) => first_stage_im_out(711),
            data_im_out(12) => first_stage_im_out(775),
            data_im_out(13) => first_stage_im_out(839),
            data_im_out(14) => first_stage_im_out(903),
            data_im_out(15) => first_stage_im_out(967),
            data_im_out(16) => first_stage_im_out(1031),
            data_im_out(17) => first_stage_im_out(1095),
            data_im_out(18) => first_stage_im_out(1159),
            data_im_out(19) => first_stage_im_out(1223),
            data_im_out(20) => first_stage_im_out(1287),
            data_im_out(21) => first_stage_im_out(1351),
            data_im_out(22) => first_stage_im_out(1415),
            data_im_out(23) => first_stage_im_out(1479),
            data_im_out(24) => first_stage_im_out(1543),
            data_im_out(25) => first_stage_im_out(1607),
            data_im_out(26) => first_stage_im_out(1671),
            data_im_out(27) => first_stage_im_out(1735),
            data_im_out(28) => first_stage_im_out(1799),
            data_im_out(29) => first_stage_im_out(1863),
            data_im_out(30) => first_stage_im_out(1927),
            data_im_out(31) => first_stage_im_out(1991)
        );

    ULFFT_PT32_8 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(8),
            data_re_in(1) => data_re_in(72),
            data_re_in(2) => data_re_in(136),
            data_re_in(3) => data_re_in(200),
            data_re_in(4) => data_re_in(264),
            data_re_in(5) => data_re_in(328),
            data_re_in(6) => data_re_in(392),
            data_re_in(7) => data_re_in(456),
            data_re_in(8) => data_re_in(520),
            data_re_in(9) => data_re_in(584),
            data_re_in(10) => data_re_in(648),
            data_re_in(11) => data_re_in(712),
            data_re_in(12) => data_re_in(776),
            data_re_in(13) => data_re_in(840),
            data_re_in(14) => data_re_in(904),
            data_re_in(15) => data_re_in(968),
            data_re_in(16) => data_re_in(1032),
            data_re_in(17) => data_re_in(1096),
            data_re_in(18) => data_re_in(1160),
            data_re_in(19) => data_re_in(1224),
            data_re_in(20) => data_re_in(1288),
            data_re_in(21) => data_re_in(1352),
            data_re_in(22) => data_re_in(1416),
            data_re_in(23) => data_re_in(1480),
            data_re_in(24) => data_re_in(1544),
            data_re_in(25) => data_re_in(1608),
            data_re_in(26) => data_re_in(1672),
            data_re_in(27) => data_re_in(1736),
            data_re_in(28) => data_re_in(1800),
            data_re_in(29) => data_re_in(1864),
            data_re_in(30) => data_re_in(1928),
            data_re_in(31) => data_re_in(1992),
            data_im_in(0) => data_im_in(8),
            data_im_in(1) => data_im_in(72),
            data_im_in(2) => data_im_in(136),
            data_im_in(3) => data_im_in(200),
            data_im_in(4) => data_im_in(264),
            data_im_in(5) => data_im_in(328),
            data_im_in(6) => data_im_in(392),
            data_im_in(7) => data_im_in(456),
            data_im_in(8) => data_im_in(520),
            data_im_in(9) => data_im_in(584),
            data_im_in(10) => data_im_in(648),
            data_im_in(11) => data_im_in(712),
            data_im_in(12) => data_im_in(776),
            data_im_in(13) => data_im_in(840),
            data_im_in(14) => data_im_in(904),
            data_im_in(15) => data_im_in(968),
            data_im_in(16) => data_im_in(1032),
            data_im_in(17) => data_im_in(1096),
            data_im_in(18) => data_im_in(1160),
            data_im_in(19) => data_im_in(1224),
            data_im_in(20) => data_im_in(1288),
            data_im_in(21) => data_im_in(1352),
            data_im_in(22) => data_im_in(1416),
            data_im_in(23) => data_im_in(1480),
            data_im_in(24) => data_im_in(1544),
            data_im_in(25) => data_im_in(1608),
            data_im_in(26) => data_im_in(1672),
            data_im_in(27) => data_im_in(1736),
            data_im_in(28) => data_im_in(1800),
            data_im_in(29) => data_im_in(1864),
            data_im_in(30) => data_im_in(1928),
            data_im_in(31) => data_im_in(1992),
            data_re_out(0) => first_stage_re_out(8),
            data_re_out(1) => first_stage_re_out(72),
            data_re_out(2) => first_stage_re_out(136),
            data_re_out(3) => first_stage_re_out(200),
            data_re_out(4) => first_stage_re_out(264),
            data_re_out(5) => first_stage_re_out(328),
            data_re_out(6) => first_stage_re_out(392),
            data_re_out(7) => first_stage_re_out(456),
            data_re_out(8) => first_stage_re_out(520),
            data_re_out(9) => first_stage_re_out(584),
            data_re_out(10) => first_stage_re_out(648),
            data_re_out(11) => first_stage_re_out(712),
            data_re_out(12) => first_stage_re_out(776),
            data_re_out(13) => first_stage_re_out(840),
            data_re_out(14) => first_stage_re_out(904),
            data_re_out(15) => first_stage_re_out(968),
            data_re_out(16) => first_stage_re_out(1032),
            data_re_out(17) => first_stage_re_out(1096),
            data_re_out(18) => first_stage_re_out(1160),
            data_re_out(19) => first_stage_re_out(1224),
            data_re_out(20) => first_stage_re_out(1288),
            data_re_out(21) => first_stage_re_out(1352),
            data_re_out(22) => first_stage_re_out(1416),
            data_re_out(23) => first_stage_re_out(1480),
            data_re_out(24) => first_stage_re_out(1544),
            data_re_out(25) => first_stage_re_out(1608),
            data_re_out(26) => first_stage_re_out(1672),
            data_re_out(27) => first_stage_re_out(1736),
            data_re_out(28) => first_stage_re_out(1800),
            data_re_out(29) => first_stage_re_out(1864),
            data_re_out(30) => first_stage_re_out(1928),
            data_re_out(31) => first_stage_re_out(1992),
            data_im_out(0) => first_stage_im_out(8),
            data_im_out(1) => first_stage_im_out(72),
            data_im_out(2) => first_stage_im_out(136),
            data_im_out(3) => first_stage_im_out(200),
            data_im_out(4) => first_stage_im_out(264),
            data_im_out(5) => first_stage_im_out(328),
            data_im_out(6) => first_stage_im_out(392),
            data_im_out(7) => first_stage_im_out(456),
            data_im_out(8) => first_stage_im_out(520),
            data_im_out(9) => first_stage_im_out(584),
            data_im_out(10) => first_stage_im_out(648),
            data_im_out(11) => first_stage_im_out(712),
            data_im_out(12) => first_stage_im_out(776),
            data_im_out(13) => first_stage_im_out(840),
            data_im_out(14) => first_stage_im_out(904),
            data_im_out(15) => first_stage_im_out(968),
            data_im_out(16) => first_stage_im_out(1032),
            data_im_out(17) => first_stage_im_out(1096),
            data_im_out(18) => first_stage_im_out(1160),
            data_im_out(19) => first_stage_im_out(1224),
            data_im_out(20) => first_stage_im_out(1288),
            data_im_out(21) => first_stage_im_out(1352),
            data_im_out(22) => first_stage_im_out(1416),
            data_im_out(23) => first_stage_im_out(1480),
            data_im_out(24) => first_stage_im_out(1544),
            data_im_out(25) => first_stage_im_out(1608),
            data_im_out(26) => first_stage_im_out(1672),
            data_im_out(27) => first_stage_im_out(1736),
            data_im_out(28) => first_stage_im_out(1800),
            data_im_out(29) => first_stage_im_out(1864),
            data_im_out(30) => first_stage_im_out(1928),
            data_im_out(31) => first_stage_im_out(1992)
        );

    ULFFT_PT32_9 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(9),
            data_re_in(1) => data_re_in(73),
            data_re_in(2) => data_re_in(137),
            data_re_in(3) => data_re_in(201),
            data_re_in(4) => data_re_in(265),
            data_re_in(5) => data_re_in(329),
            data_re_in(6) => data_re_in(393),
            data_re_in(7) => data_re_in(457),
            data_re_in(8) => data_re_in(521),
            data_re_in(9) => data_re_in(585),
            data_re_in(10) => data_re_in(649),
            data_re_in(11) => data_re_in(713),
            data_re_in(12) => data_re_in(777),
            data_re_in(13) => data_re_in(841),
            data_re_in(14) => data_re_in(905),
            data_re_in(15) => data_re_in(969),
            data_re_in(16) => data_re_in(1033),
            data_re_in(17) => data_re_in(1097),
            data_re_in(18) => data_re_in(1161),
            data_re_in(19) => data_re_in(1225),
            data_re_in(20) => data_re_in(1289),
            data_re_in(21) => data_re_in(1353),
            data_re_in(22) => data_re_in(1417),
            data_re_in(23) => data_re_in(1481),
            data_re_in(24) => data_re_in(1545),
            data_re_in(25) => data_re_in(1609),
            data_re_in(26) => data_re_in(1673),
            data_re_in(27) => data_re_in(1737),
            data_re_in(28) => data_re_in(1801),
            data_re_in(29) => data_re_in(1865),
            data_re_in(30) => data_re_in(1929),
            data_re_in(31) => data_re_in(1993),
            data_im_in(0) => data_im_in(9),
            data_im_in(1) => data_im_in(73),
            data_im_in(2) => data_im_in(137),
            data_im_in(3) => data_im_in(201),
            data_im_in(4) => data_im_in(265),
            data_im_in(5) => data_im_in(329),
            data_im_in(6) => data_im_in(393),
            data_im_in(7) => data_im_in(457),
            data_im_in(8) => data_im_in(521),
            data_im_in(9) => data_im_in(585),
            data_im_in(10) => data_im_in(649),
            data_im_in(11) => data_im_in(713),
            data_im_in(12) => data_im_in(777),
            data_im_in(13) => data_im_in(841),
            data_im_in(14) => data_im_in(905),
            data_im_in(15) => data_im_in(969),
            data_im_in(16) => data_im_in(1033),
            data_im_in(17) => data_im_in(1097),
            data_im_in(18) => data_im_in(1161),
            data_im_in(19) => data_im_in(1225),
            data_im_in(20) => data_im_in(1289),
            data_im_in(21) => data_im_in(1353),
            data_im_in(22) => data_im_in(1417),
            data_im_in(23) => data_im_in(1481),
            data_im_in(24) => data_im_in(1545),
            data_im_in(25) => data_im_in(1609),
            data_im_in(26) => data_im_in(1673),
            data_im_in(27) => data_im_in(1737),
            data_im_in(28) => data_im_in(1801),
            data_im_in(29) => data_im_in(1865),
            data_im_in(30) => data_im_in(1929),
            data_im_in(31) => data_im_in(1993),
            data_re_out(0) => first_stage_re_out(9),
            data_re_out(1) => first_stage_re_out(73),
            data_re_out(2) => first_stage_re_out(137),
            data_re_out(3) => first_stage_re_out(201),
            data_re_out(4) => first_stage_re_out(265),
            data_re_out(5) => first_stage_re_out(329),
            data_re_out(6) => first_stage_re_out(393),
            data_re_out(7) => first_stage_re_out(457),
            data_re_out(8) => first_stage_re_out(521),
            data_re_out(9) => first_stage_re_out(585),
            data_re_out(10) => first_stage_re_out(649),
            data_re_out(11) => first_stage_re_out(713),
            data_re_out(12) => first_stage_re_out(777),
            data_re_out(13) => first_stage_re_out(841),
            data_re_out(14) => first_stage_re_out(905),
            data_re_out(15) => first_stage_re_out(969),
            data_re_out(16) => first_stage_re_out(1033),
            data_re_out(17) => first_stage_re_out(1097),
            data_re_out(18) => first_stage_re_out(1161),
            data_re_out(19) => first_stage_re_out(1225),
            data_re_out(20) => first_stage_re_out(1289),
            data_re_out(21) => first_stage_re_out(1353),
            data_re_out(22) => first_stage_re_out(1417),
            data_re_out(23) => first_stage_re_out(1481),
            data_re_out(24) => first_stage_re_out(1545),
            data_re_out(25) => first_stage_re_out(1609),
            data_re_out(26) => first_stage_re_out(1673),
            data_re_out(27) => first_stage_re_out(1737),
            data_re_out(28) => first_stage_re_out(1801),
            data_re_out(29) => first_stage_re_out(1865),
            data_re_out(30) => first_stage_re_out(1929),
            data_re_out(31) => first_stage_re_out(1993),
            data_im_out(0) => first_stage_im_out(9),
            data_im_out(1) => first_stage_im_out(73),
            data_im_out(2) => first_stage_im_out(137),
            data_im_out(3) => first_stage_im_out(201),
            data_im_out(4) => first_stage_im_out(265),
            data_im_out(5) => first_stage_im_out(329),
            data_im_out(6) => first_stage_im_out(393),
            data_im_out(7) => first_stage_im_out(457),
            data_im_out(8) => first_stage_im_out(521),
            data_im_out(9) => first_stage_im_out(585),
            data_im_out(10) => first_stage_im_out(649),
            data_im_out(11) => first_stage_im_out(713),
            data_im_out(12) => first_stage_im_out(777),
            data_im_out(13) => first_stage_im_out(841),
            data_im_out(14) => first_stage_im_out(905),
            data_im_out(15) => first_stage_im_out(969),
            data_im_out(16) => first_stage_im_out(1033),
            data_im_out(17) => first_stage_im_out(1097),
            data_im_out(18) => first_stage_im_out(1161),
            data_im_out(19) => first_stage_im_out(1225),
            data_im_out(20) => first_stage_im_out(1289),
            data_im_out(21) => first_stage_im_out(1353),
            data_im_out(22) => first_stage_im_out(1417),
            data_im_out(23) => first_stage_im_out(1481),
            data_im_out(24) => first_stage_im_out(1545),
            data_im_out(25) => first_stage_im_out(1609),
            data_im_out(26) => first_stage_im_out(1673),
            data_im_out(27) => first_stage_im_out(1737),
            data_im_out(28) => first_stage_im_out(1801),
            data_im_out(29) => first_stage_im_out(1865),
            data_im_out(30) => first_stage_im_out(1929),
            data_im_out(31) => first_stage_im_out(1993)
        );

    ULFFT_PT32_10 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(10),
            data_re_in(1) => data_re_in(74),
            data_re_in(2) => data_re_in(138),
            data_re_in(3) => data_re_in(202),
            data_re_in(4) => data_re_in(266),
            data_re_in(5) => data_re_in(330),
            data_re_in(6) => data_re_in(394),
            data_re_in(7) => data_re_in(458),
            data_re_in(8) => data_re_in(522),
            data_re_in(9) => data_re_in(586),
            data_re_in(10) => data_re_in(650),
            data_re_in(11) => data_re_in(714),
            data_re_in(12) => data_re_in(778),
            data_re_in(13) => data_re_in(842),
            data_re_in(14) => data_re_in(906),
            data_re_in(15) => data_re_in(970),
            data_re_in(16) => data_re_in(1034),
            data_re_in(17) => data_re_in(1098),
            data_re_in(18) => data_re_in(1162),
            data_re_in(19) => data_re_in(1226),
            data_re_in(20) => data_re_in(1290),
            data_re_in(21) => data_re_in(1354),
            data_re_in(22) => data_re_in(1418),
            data_re_in(23) => data_re_in(1482),
            data_re_in(24) => data_re_in(1546),
            data_re_in(25) => data_re_in(1610),
            data_re_in(26) => data_re_in(1674),
            data_re_in(27) => data_re_in(1738),
            data_re_in(28) => data_re_in(1802),
            data_re_in(29) => data_re_in(1866),
            data_re_in(30) => data_re_in(1930),
            data_re_in(31) => data_re_in(1994),
            data_im_in(0) => data_im_in(10),
            data_im_in(1) => data_im_in(74),
            data_im_in(2) => data_im_in(138),
            data_im_in(3) => data_im_in(202),
            data_im_in(4) => data_im_in(266),
            data_im_in(5) => data_im_in(330),
            data_im_in(6) => data_im_in(394),
            data_im_in(7) => data_im_in(458),
            data_im_in(8) => data_im_in(522),
            data_im_in(9) => data_im_in(586),
            data_im_in(10) => data_im_in(650),
            data_im_in(11) => data_im_in(714),
            data_im_in(12) => data_im_in(778),
            data_im_in(13) => data_im_in(842),
            data_im_in(14) => data_im_in(906),
            data_im_in(15) => data_im_in(970),
            data_im_in(16) => data_im_in(1034),
            data_im_in(17) => data_im_in(1098),
            data_im_in(18) => data_im_in(1162),
            data_im_in(19) => data_im_in(1226),
            data_im_in(20) => data_im_in(1290),
            data_im_in(21) => data_im_in(1354),
            data_im_in(22) => data_im_in(1418),
            data_im_in(23) => data_im_in(1482),
            data_im_in(24) => data_im_in(1546),
            data_im_in(25) => data_im_in(1610),
            data_im_in(26) => data_im_in(1674),
            data_im_in(27) => data_im_in(1738),
            data_im_in(28) => data_im_in(1802),
            data_im_in(29) => data_im_in(1866),
            data_im_in(30) => data_im_in(1930),
            data_im_in(31) => data_im_in(1994),
            data_re_out(0) => first_stage_re_out(10),
            data_re_out(1) => first_stage_re_out(74),
            data_re_out(2) => first_stage_re_out(138),
            data_re_out(3) => first_stage_re_out(202),
            data_re_out(4) => first_stage_re_out(266),
            data_re_out(5) => first_stage_re_out(330),
            data_re_out(6) => first_stage_re_out(394),
            data_re_out(7) => first_stage_re_out(458),
            data_re_out(8) => first_stage_re_out(522),
            data_re_out(9) => first_stage_re_out(586),
            data_re_out(10) => first_stage_re_out(650),
            data_re_out(11) => first_stage_re_out(714),
            data_re_out(12) => first_stage_re_out(778),
            data_re_out(13) => first_stage_re_out(842),
            data_re_out(14) => first_stage_re_out(906),
            data_re_out(15) => first_stage_re_out(970),
            data_re_out(16) => first_stage_re_out(1034),
            data_re_out(17) => first_stage_re_out(1098),
            data_re_out(18) => first_stage_re_out(1162),
            data_re_out(19) => first_stage_re_out(1226),
            data_re_out(20) => first_stage_re_out(1290),
            data_re_out(21) => first_stage_re_out(1354),
            data_re_out(22) => first_stage_re_out(1418),
            data_re_out(23) => first_stage_re_out(1482),
            data_re_out(24) => first_stage_re_out(1546),
            data_re_out(25) => first_stage_re_out(1610),
            data_re_out(26) => first_stage_re_out(1674),
            data_re_out(27) => first_stage_re_out(1738),
            data_re_out(28) => first_stage_re_out(1802),
            data_re_out(29) => first_stage_re_out(1866),
            data_re_out(30) => first_stage_re_out(1930),
            data_re_out(31) => first_stage_re_out(1994),
            data_im_out(0) => first_stage_im_out(10),
            data_im_out(1) => first_stage_im_out(74),
            data_im_out(2) => first_stage_im_out(138),
            data_im_out(3) => first_stage_im_out(202),
            data_im_out(4) => first_stage_im_out(266),
            data_im_out(5) => first_stage_im_out(330),
            data_im_out(6) => first_stage_im_out(394),
            data_im_out(7) => first_stage_im_out(458),
            data_im_out(8) => first_stage_im_out(522),
            data_im_out(9) => first_stage_im_out(586),
            data_im_out(10) => first_stage_im_out(650),
            data_im_out(11) => first_stage_im_out(714),
            data_im_out(12) => first_stage_im_out(778),
            data_im_out(13) => first_stage_im_out(842),
            data_im_out(14) => first_stage_im_out(906),
            data_im_out(15) => first_stage_im_out(970),
            data_im_out(16) => first_stage_im_out(1034),
            data_im_out(17) => first_stage_im_out(1098),
            data_im_out(18) => first_stage_im_out(1162),
            data_im_out(19) => first_stage_im_out(1226),
            data_im_out(20) => first_stage_im_out(1290),
            data_im_out(21) => first_stage_im_out(1354),
            data_im_out(22) => first_stage_im_out(1418),
            data_im_out(23) => first_stage_im_out(1482),
            data_im_out(24) => first_stage_im_out(1546),
            data_im_out(25) => first_stage_im_out(1610),
            data_im_out(26) => first_stage_im_out(1674),
            data_im_out(27) => first_stage_im_out(1738),
            data_im_out(28) => first_stage_im_out(1802),
            data_im_out(29) => first_stage_im_out(1866),
            data_im_out(30) => first_stage_im_out(1930),
            data_im_out(31) => first_stage_im_out(1994)
        );

    ULFFT_PT32_11 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(11),
            data_re_in(1) => data_re_in(75),
            data_re_in(2) => data_re_in(139),
            data_re_in(3) => data_re_in(203),
            data_re_in(4) => data_re_in(267),
            data_re_in(5) => data_re_in(331),
            data_re_in(6) => data_re_in(395),
            data_re_in(7) => data_re_in(459),
            data_re_in(8) => data_re_in(523),
            data_re_in(9) => data_re_in(587),
            data_re_in(10) => data_re_in(651),
            data_re_in(11) => data_re_in(715),
            data_re_in(12) => data_re_in(779),
            data_re_in(13) => data_re_in(843),
            data_re_in(14) => data_re_in(907),
            data_re_in(15) => data_re_in(971),
            data_re_in(16) => data_re_in(1035),
            data_re_in(17) => data_re_in(1099),
            data_re_in(18) => data_re_in(1163),
            data_re_in(19) => data_re_in(1227),
            data_re_in(20) => data_re_in(1291),
            data_re_in(21) => data_re_in(1355),
            data_re_in(22) => data_re_in(1419),
            data_re_in(23) => data_re_in(1483),
            data_re_in(24) => data_re_in(1547),
            data_re_in(25) => data_re_in(1611),
            data_re_in(26) => data_re_in(1675),
            data_re_in(27) => data_re_in(1739),
            data_re_in(28) => data_re_in(1803),
            data_re_in(29) => data_re_in(1867),
            data_re_in(30) => data_re_in(1931),
            data_re_in(31) => data_re_in(1995),
            data_im_in(0) => data_im_in(11),
            data_im_in(1) => data_im_in(75),
            data_im_in(2) => data_im_in(139),
            data_im_in(3) => data_im_in(203),
            data_im_in(4) => data_im_in(267),
            data_im_in(5) => data_im_in(331),
            data_im_in(6) => data_im_in(395),
            data_im_in(7) => data_im_in(459),
            data_im_in(8) => data_im_in(523),
            data_im_in(9) => data_im_in(587),
            data_im_in(10) => data_im_in(651),
            data_im_in(11) => data_im_in(715),
            data_im_in(12) => data_im_in(779),
            data_im_in(13) => data_im_in(843),
            data_im_in(14) => data_im_in(907),
            data_im_in(15) => data_im_in(971),
            data_im_in(16) => data_im_in(1035),
            data_im_in(17) => data_im_in(1099),
            data_im_in(18) => data_im_in(1163),
            data_im_in(19) => data_im_in(1227),
            data_im_in(20) => data_im_in(1291),
            data_im_in(21) => data_im_in(1355),
            data_im_in(22) => data_im_in(1419),
            data_im_in(23) => data_im_in(1483),
            data_im_in(24) => data_im_in(1547),
            data_im_in(25) => data_im_in(1611),
            data_im_in(26) => data_im_in(1675),
            data_im_in(27) => data_im_in(1739),
            data_im_in(28) => data_im_in(1803),
            data_im_in(29) => data_im_in(1867),
            data_im_in(30) => data_im_in(1931),
            data_im_in(31) => data_im_in(1995),
            data_re_out(0) => first_stage_re_out(11),
            data_re_out(1) => first_stage_re_out(75),
            data_re_out(2) => first_stage_re_out(139),
            data_re_out(3) => first_stage_re_out(203),
            data_re_out(4) => first_stage_re_out(267),
            data_re_out(5) => first_stage_re_out(331),
            data_re_out(6) => first_stage_re_out(395),
            data_re_out(7) => first_stage_re_out(459),
            data_re_out(8) => first_stage_re_out(523),
            data_re_out(9) => first_stage_re_out(587),
            data_re_out(10) => first_stage_re_out(651),
            data_re_out(11) => first_stage_re_out(715),
            data_re_out(12) => first_stage_re_out(779),
            data_re_out(13) => first_stage_re_out(843),
            data_re_out(14) => first_stage_re_out(907),
            data_re_out(15) => first_stage_re_out(971),
            data_re_out(16) => first_stage_re_out(1035),
            data_re_out(17) => first_stage_re_out(1099),
            data_re_out(18) => first_stage_re_out(1163),
            data_re_out(19) => first_stage_re_out(1227),
            data_re_out(20) => first_stage_re_out(1291),
            data_re_out(21) => first_stage_re_out(1355),
            data_re_out(22) => first_stage_re_out(1419),
            data_re_out(23) => first_stage_re_out(1483),
            data_re_out(24) => first_stage_re_out(1547),
            data_re_out(25) => first_stage_re_out(1611),
            data_re_out(26) => first_stage_re_out(1675),
            data_re_out(27) => first_stage_re_out(1739),
            data_re_out(28) => first_stage_re_out(1803),
            data_re_out(29) => first_stage_re_out(1867),
            data_re_out(30) => first_stage_re_out(1931),
            data_re_out(31) => first_stage_re_out(1995),
            data_im_out(0) => first_stage_im_out(11),
            data_im_out(1) => first_stage_im_out(75),
            data_im_out(2) => first_stage_im_out(139),
            data_im_out(3) => first_stage_im_out(203),
            data_im_out(4) => first_stage_im_out(267),
            data_im_out(5) => first_stage_im_out(331),
            data_im_out(6) => first_stage_im_out(395),
            data_im_out(7) => first_stage_im_out(459),
            data_im_out(8) => first_stage_im_out(523),
            data_im_out(9) => first_stage_im_out(587),
            data_im_out(10) => first_stage_im_out(651),
            data_im_out(11) => first_stage_im_out(715),
            data_im_out(12) => first_stage_im_out(779),
            data_im_out(13) => first_stage_im_out(843),
            data_im_out(14) => first_stage_im_out(907),
            data_im_out(15) => first_stage_im_out(971),
            data_im_out(16) => first_stage_im_out(1035),
            data_im_out(17) => first_stage_im_out(1099),
            data_im_out(18) => first_stage_im_out(1163),
            data_im_out(19) => first_stage_im_out(1227),
            data_im_out(20) => first_stage_im_out(1291),
            data_im_out(21) => first_stage_im_out(1355),
            data_im_out(22) => first_stage_im_out(1419),
            data_im_out(23) => first_stage_im_out(1483),
            data_im_out(24) => first_stage_im_out(1547),
            data_im_out(25) => first_stage_im_out(1611),
            data_im_out(26) => first_stage_im_out(1675),
            data_im_out(27) => first_stage_im_out(1739),
            data_im_out(28) => first_stage_im_out(1803),
            data_im_out(29) => first_stage_im_out(1867),
            data_im_out(30) => first_stage_im_out(1931),
            data_im_out(31) => first_stage_im_out(1995)
        );

    ULFFT_PT32_12 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(12),
            data_re_in(1) => data_re_in(76),
            data_re_in(2) => data_re_in(140),
            data_re_in(3) => data_re_in(204),
            data_re_in(4) => data_re_in(268),
            data_re_in(5) => data_re_in(332),
            data_re_in(6) => data_re_in(396),
            data_re_in(7) => data_re_in(460),
            data_re_in(8) => data_re_in(524),
            data_re_in(9) => data_re_in(588),
            data_re_in(10) => data_re_in(652),
            data_re_in(11) => data_re_in(716),
            data_re_in(12) => data_re_in(780),
            data_re_in(13) => data_re_in(844),
            data_re_in(14) => data_re_in(908),
            data_re_in(15) => data_re_in(972),
            data_re_in(16) => data_re_in(1036),
            data_re_in(17) => data_re_in(1100),
            data_re_in(18) => data_re_in(1164),
            data_re_in(19) => data_re_in(1228),
            data_re_in(20) => data_re_in(1292),
            data_re_in(21) => data_re_in(1356),
            data_re_in(22) => data_re_in(1420),
            data_re_in(23) => data_re_in(1484),
            data_re_in(24) => data_re_in(1548),
            data_re_in(25) => data_re_in(1612),
            data_re_in(26) => data_re_in(1676),
            data_re_in(27) => data_re_in(1740),
            data_re_in(28) => data_re_in(1804),
            data_re_in(29) => data_re_in(1868),
            data_re_in(30) => data_re_in(1932),
            data_re_in(31) => data_re_in(1996),
            data_im_in(0) => data_im_in(12),
            data_im_in(1) => data_im_in(76),
            data_im_in(2) => data_im_in(140),
            data_im_in(3) => data_im_in(204),
            data_im_in(4) => data_im_in(268),
            data_im_in(5) => data_im_in(332),
            data_im_in(6) => data_im_in(396),
            data_im_in(7) => data_im_in(460),
            data_im_in(8) => data_im_in(524),
            data_im_in(9) => data_im_in(588),
            data_im_in(10) => data_im_in(652),
            data_im_in(11) => data_im_in(716),
            data_im_in(12) => data_im_in(780),
            data_im_in(13) => data_im_in(844),
            data_im_in(14) => data_im_in(908),
            data_im_in(15) => data_im_in(972),
            data_im_in(16) => data_im_in(1036),
            data_im_in(17) => data_im_in(1100),
            data_im_in(18) => data_im_in(1164),
            data_im_in(19) => data_im_in(1228),
            data_im_in(20) => data_im_in(1292),
            data_im_in(21) => data_im_in(1356),
            data_im_in(22) => data_im_in(1420),
            data_im_in(23) => data_im_in(1484),
            data_im_in(24) => data_im_in(1548),
            data_im_in(25) => data_im_in(1612),
            data_im_in(26) => data_im_in(1676),
            data_im_in(27) => data_im_in(1740),
            data_im_in(28) => data_im_in(1804),
            data_im_in(29) => data_im_in(1868),
            data_im_in(30) => data_im_in(1932),
            data_im_in(31) => data_im_in(1996),
            data_re_out(0) => first_stage_re_out(12),
            data_re_out(1) => first_stage_re_out(76),
            data_re_out(2) => first_stage_re_out(140),
            data_re_out(3) => first_stage_re_out(204),
            data_re_out(4) => first_stage_re_out(268),
            data_re_out(5) => first_stage_re_out(332),
            data_re_out(6) => first_stage_re_out(396),
            data_re_out(7) => first_stage_re_out(460),
            data_re_out(8) => first_stage_re_out(524),
            data_re_out(9) => first_stage_re_out(588),
            data_re_out(10) => first_stage_re_out(652),
            data_re_out(11) => first_stage_re_out(716),
            data_re_out(12) => first_stage_re_out(780),
            data_re_out(13) => first_stage_re_out(844),
            data_re_out(14) => first_stage_re_out(908),
            data_re_out(15) => first_stage_re_out(972),
            data_re_out(16) => first_stage_re_out(1036),
            data_re_out(17) => first_stage_re_out(1100),
            data_re_out(18) => first_stage_re_out(1164),
            data_re_out(19) => first_stage_re_out(1228),
            data_re_out(20) => first_stage_re_out(1292),
            data_re_out(21) => first_stage_re_out(1356),
            data_re_out(22) => first_stage_re_out(1420),
            data_re_out(23) => first_stage_re_out(1484),
            data_re_out(24) => first_stage_re_out(1548),
            data_re_out(25) => first_stage_re_out(1612),
            data_re_out(26) => first_stage_re_out(1676),
            data_re_out(27) => first_stage_re_out(1740),
            data_re_out(28) => first_stage_re_out(1804),
            data_re_out(29) => first_stage_re_out(1868),
            data_re_out(30) => first_stage_re_out(1932),
            data_re_out(31) => first_stage_re_out(1996),
            data_im_out(0) => first_stage_im_out(12),
            data_im_out(1) => first_stage_im_out(76),
            data_im_out(2) => first_stage_im_out(140),
            data_im_out(3) => first_stage_im_out(204),
            data_im_out(4) => first_stage_im_out(268),
            data_im_out(5) => first_stage_im_out(332),
            data_im_out(6) => first_stage_im_out(396),
            data_im_out(7) => first_stage_im_out(460),
            data_im_out(8) => first_stage_im_out(524),
            data_im_out(9) => first_stage_im_out(588),
            data_im_out(10) => first_stage_im_out(652),
            data_im_out(11) => first_stage_im_out(716),
            data_im_out(12) => first_stage_im_out(780),
            data_im_out(13) => first_stage_im_out(844),
            data_im_out(14) => first_stage_im_out(908),
            data_im_out(15) => first_stage_im_out(972),
            data_im_out(16) => first_stage_im_out(1036),
            data_im_out(17) => first_stage_im_out(1100),
            data_im_out(18) => first_stage_im_out(1164),
            data_im_out(19) => first_stage_im_out(1228),
            data_im_out(20) => first_stage_im_out(1292),
            data_im_out(21) => first_stage_im_out(1356),
            data_im_out(22) => first_stage_im_out(1420),
            data_im_out(23) => first_stage_im_out(1484),
            data_im_out(24) => first_stage_im_out(1548),
            data_im_out(25) => first_stage_im_out(1612),
            data_im_out(26) => first_stage_im_out(1676),
            data_im_out(27) => first_stage_im_out(1740),
            data_im_out(28) => first_stage_im_out(1804),
            data_im_out(29) => first_stage_im_out(1868),
            data_im_out(30) => first_stage_im_out(1932),
            data_im_out(31) => first_stage_im_out(1996)
        );

    ULFFT_PT32_13 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(13),
            data_re_in(1) => data_re_in(77),
            data_re_in(2) => data_re_in(141),
            data_re_in(3) => data_re_in(205),
            data_re_in(4) => data_re_in(269),
            data_re_in(5) => data_re_in(333),
            data_re_in(6) => data_re_in(397),
            data_re_in(7) => data_re_in(461),
            data_re_in(8) => data_re_in(525),
            data_re_in(9) => data_re_in(589),
            data_re_in(10) => data_re_in(653),
            data_re_in(11) => data_re_in(717),
            data_re_in(12) => data_re_in(781),
            data_re_in(13) => data_re_in(845),
            data_re_in(14) => data_re_in(909),
            data_re_in(15) => data_re_in(973),
            data_re_in(16) => data_re_in(1037),
            data_re_in(17) => data_re_in(1101),
            data_re_in(18) => data_re_in(1165),
            data_re_in(19) => data_re_in(1229),
            data_re_in(20) => data_re_in(1293),
            data_re_in(21) => data_re_in(1357),
            data_re_in(22) => data_re_in(1421),
            data_re_in(23) => data_re_in(1485),
            data_re_in(24) => data_re_in(1549),
            data_re_in(25) => data_re_in(1613),
            data_re_in(26) => data_re_in(1677),
            data_re_in(27) => data_re_in(1741),
            data_re_in(28) => data_re_in(1805),
            data_re_in(29) => data_re_in(1869),
            data_re_in(30) => data_re_in(1933),
            data_re_in(31) => data_re_in(1997),
            data_im_in(0) => data_im_in(13),
            data_im_in(1) => data_im_in(77),
            data_im_in(2) => data_im_in(141),
            data_im_in(3) => data_im_in(205),
            data_im_in(4) => data_im_in(269),
            data_im_in(5) => data_im_in(333),
            data_im_in(6) => data_im_in(397),
            data_im_in(7) => data_im_in(461),
            data_im_in(8) => data_im_in(525),
            data_im_in(9) => data_im_in(589),
            data_im_in(10) => data_im_in(653),
            data_im_in(11) => data_im_in(717),
            data_im_in(12) => data_im_in(781),
            data_im_in(13) => data_im_in(845),
            data_im_in(14) => data_im_in(909),
            data_im_in(15) => data_im_in(973),
            data_im_in(16) => data_im_in(1037),
            data_im_in(17) => data_im_in(1101),
            data_im_in(18) => data_im_in(1165),
            data_im_in(19) => data_im_in(1229),
            data_im_in(20) => data_im_in(1293),
            data_im_in(21) => data_im_in(1357),
            data_im_in(22) => data_im_in(1421),
            data_im_in(23) => data_im_in(1485),
            data_im_in(24) => data_im_in(1549),
            data_im_in(25) => data_im_in(1613),
            data_im_in(26) => data_im_in(1677),
            data_im_in(27) => data_im_in(1741),
            data_im_in(28) => data_im_in(1805),
            data_im_in(29) => data_im_in(1869),
            data_im_in(30) => data_im_in(1933),
            data_im_in(31) => data_im_in(1997),
            data_re_out(0) => first_stage_re_out(13),
            data_re_out(1) => first_stage_re_out(77),
            data_re_out(2) => first_stage_re_out(141),
            data_re_out(3) => first_stage_re_out(205),
            data_re_out(4) => first_stage_re_out(269),
            data_re_out(5) => first_stage_re_out(333),
            data_re_out(6) => first_stage_re_out(397),
            data_re_out(7) => first_stage_re_out(461),
            data_re_out(8) => first_stage_re_out(525),
            data_re_out(9) => first_stage_re_out(589),
            data_re_out(10) => first_stage_re_out(653),
            data_re_out(11) => first_stage_re_out(717),
            data_re_out(12) => first_stage_re_out(781),
            data_re_out(13) => first_stage_re_out(845),
            data_re_out(14) => first_stage_re_out(909),
            data_re_out(15) => first_stage_re_out(973),
            data_re_out(16) => first_stage_re_out(1037),
            data_re_out(17) => first_stage_re_out(1101),
            data_re_out(18) => first_stage_re_out(1165),
            data_re_out(19) => first_stage_re_out(1229),
            data_re_out(20) => first_stage_re_out(1293),
            data_re_out(21) => first_stage_re_out(1357),
            data_re_out(22) => first_stage_re_out(1421),
            data_re_out(23) => first_stage_re_out(1485),
            data_re_out(24) => first_stage_re_out(1549),
            data_re_out(25) => first_stage_re_out(1613),
            data_re_out(26) => first_stage_re_out(1677),
            data_re_out(27) => first_stage_re_out(1741),
            data_re_out(28) => first_stage_re_out(1805),
            data_re_out(29) => first_stage_re_out(1869),
            data_re_out(30) => first_stage_re_out(1933),
            data_re_out(31) => first_stage_re_out(1997),
            data_im_out(0) => first_stage_im_out(13),
            data_im_out(1) => first_stage_im_out(77),
            data_im_out(2) => first_stage_im_out(141),
            data_im_out(3) => first_stage_im_out(205),
            data_im_out(4) => first_stage_im_out(269),
            data_im_out(5) => first_stage_im_out(333),
            data_im_out(6) => first_stage_im_out(397),
            data_im_out(7) => first_stage_im_out(461),
            data_im_out(8) => first_stage_im_out(525),
            data_im_out(9) => first_stage_im_out(589),
            data_im_out(10) => first_stage_im_out(653),
            data_im_out(11) => first_stage_im_out(717),
            data_im_out(12) => first_stage_im_out(781),
            data_im_out(13) => first_stage_im_out(845),
            data_im_out(14) => first_stage_im_out(909),
            data_im_out(15) => first_stage_im_out(973),
            data_im_out(16) => first_stage_im_out(1037),
            data_im_out(17) => first_stage_im_out(1101),
            data_im_out(18) => first_stage_im_out(1165),
            data_im_out(19) => first_stage_im_out(1229),
            data_im_out(20) => first_stage_im_out(1293),
            data_im_out(21) => first_stage_im_out(1357),
            data_im_out(22) => first_stage_im_out(1421),
            data_im_out(23) => first_stage_im_out(1485),
            data_im_out(24) => first_stage_im_out(1549),
            data_im_out(25) => first_stage_im_out(1613),
            data_im_out(26) => first_stage_im_out(1677),
            data_im_out(27) => first_stage_im_out(1741),
            data_im_out(28) => first_stage_im_out(1805),
            data_im_out(29) => first_stage_im_out(1869),
            data_im_out(30) => first_stage_im_out(1933),
            data_im_out(31) => first_stage_im_out(1997)
        );

    ULFFT_PT32_14 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(14),
            data_re_in(1) => data_re_in(78),
            data_re_in(2) => data_re_in(142),
            data_re_in(3) => data_re_in(206),
            data_re_in(4) => data_re_in(270),
            data_re_in(5) => data_re_in(334),
            data_re_in(6) => data_re_in(398),
            data_re_in(7) => data_re_in(462),
            data_re_in(8) => data_re_in(526),
            data_re_in(9) => data_re_in(590),
            data_re_in(10) => data_re_in(654),
            data_re_in(11) => data_re_in(718),
            data_re_in(12) => data_re_in(782),
            data_re_in(13) => data_re_in(846),
            data_re_in(14) => data_re_in(910),
            data_re_in(15) => data_re_in(974),
            data_re_in(16) => data_re_in(1038),
            data_re_in(17) => data_re_in(1102),
            data_re_in(18) => data_re_in(1166),
            data_re_in(19) => data_re_in(1230),
            data_re_in(20) => data_re_in(1294),
            data_re_in(21) => data_re_in(1358),
            data_re_in(22) => data_re_in(1422),
            data_re_in(23) => data_re_in(1486),
            data_re_in(24) => data_re_in(1550),
            data_re_in(25) => data_re_in(1614),
            data_re_in(26) => data_re_in(1678),
            data_re_in(27) => data_re_in(1742),
            data_re_in(28) => data_re_in(1806),
            data_re_in(29) => data_re_in(1870),
            data_re_in(30) => data_re_in(1934),
            data_re_in(31) => data_re_in(1998),
            data_im_in(0) => data_im_in(14),
            data_im_in(1) => data_im_in(78),
            data_im_in(2) => data_im_in(142),
            data_im_in(3) => data_im_in(206),
            data_im_in(4) => data_im_in(270),
            data_im_in(5) => data_im_in(334),
            data_im_in(6) => data_im_in(398),
            data_im_in(7) => data_im_in(462),
            data_im_in(8) => data_im_in(526),
            data_im_in(9) => data_im_in(590),
            data_im_in(10) => data_im_in(654),
            data_im_in(11) => data_im_in(718),
            data_im_in(12) => data_im_in(782),
            data_im_in(13) => data_im_in(846),
            data_im_in(14) => data_im_in(910),
            data_im_in(15) => data_im_in(974),
            data_im_in(16) => data_im_in(1038),
            data_im_in(17) => data_im_in(1102),
            data_im_in(18) => data_im_in(1166),
            data_im_in(19) => data_im_in(1230),
            data_im_in(20) => data_im_in(1294),
            data_im_in(21) => data_im_in(1358),
            data_im_in(22) => data_im_in(1422),
            data_im_in(23) => data_im_in(1486),
            data_im_in(24) => data_im_in(1550),
            data_im_in(25) => data_im_in(1614),
            data_im_in(26) => data_im_in(1678),
            data_im_in(27) => data_im_in(1742),
            data_im_in(28) => data_im_in(1806),
            data_im_in(29) => data_im_in(1870),
            data_im_in(30) => data_im_in(1934),
            data_im_in(31) => data_im_in(1998),
            data_re_out(0) => first_stage_re_out(14),
            data_re_out(1) => first_stage_re_out(78),
            data_re_out(2) => first_stage_re_out(142),
            data_re_out(3) => first_stage_re_out(206),
            data_re_out(4) => first_stage_re_out(270),
            data_re_out(5) => first_stage_re_out(334),
            data_re_out(6) => first_stage_re_out(398),
            data_re_out(7) => first_stage_re_out(462),
            data_re_out(8) => first_stage_re_out(526),
            data_re_out(9) => first_stage_re_out(590),
            data_re_out(10) => first_stage_re_out(654),
            data_re_out(11) => first_stage_re_out(718),
            data_re_out(12) => first_stage_re_out(782),
            data_re_out(13) => first_stage_re_out(846),
            data_re_out(14) => first_stage_re_out(910),
            data_re_out(15) => first_stage_re_out(974),
            data_re_out(16) => first_stage_re_out(1038),
            data_re_out(17) => first_stage_re_out(1102),
            data_re_out(18) => first_stage_re_out(1166),
            data_re_out(19) => first_stage_re_out(1230),
            data_re_out(20) => first_stage_re_out(1294),
            data_re_out(21) => first_stage_re_out(1358),
            data_re_out(22) => first_stage_re_out(1422),
            data_re_out(23) => first_stage_re_out(1486),
            data_re_out(24) => first_stage_re_out(1550),
            data_re_out(25) => first_stage_re_out(1614),
            data_re_out(26) => first_stage_re_out(1678),
            data_re_out(27) => first_stage_re_out(1742),
            data_re_out(28) => first_stage_re_out(1806),
            data_re_out(29) => first_stage_re_out(1870),
            data_re_out(30) => first_stage_re_out(1934),
            data_re_out(31) => first_stage_re_out(1998),
            data_im_out(0) => first_stage_im_out(14),
            data_im_out(1) => first_stage_im_out(78),
            data_im_out(2) => first_stage_im_out(142),
            data_im_out(3) => first_stage_im_out(206),
            data_im_out(4) => first_stage_im_out(270),
            data_im_out(5) => first_stage_im_out(334),
            data_im_out(6) => first_stage_im_out(398),
            data_im_out(7) => first_stage_im_out(462),
            data_im_out(8) => first_stage_im_out(526),
            data_im_out(9) => first_stage_im_out(590),
            data_im_out(10) => first_stage_im_out(654),
            data_im_out(11) => first_stage_im_out(718),
            data_im_out(12) => first_stage_im_out(782),
            data_im_out(13) => first_stage_im_out(846),
            data_im_out(14) => first_stage_im_out(910),
            data_im_out(15) => first_stage_im_out(974),
            data_im_out(16) => first_stage_im_out(1038),
            data_im_out(17) => first_stage_im_out(1102),
            data_im_out(18) => first_stage_im_out(1166),
            data_im_out(19) => first_stage_im_out(1230),
            data_im_out(20) => first_stage_im_out(1294),
            data_im_out(21) => first_stage_im_out(1358),
            data_im_out(22) => first_stage_im_out(1422),
            data_im_out(23) => first_stage_im_out(1486),
            data_im_out(24) => first_stage_im_out(1550),
            data_im_out(25) => first_stage_im_out(1614),
            data_im_out(26) => first_stage_im_out(1678),
            data_im_out(27) => first_stage_im_out(1742),
            data_im_out(28) => first_stage_im_out(1806),
            data_im_out(29) => first_stage_im_out(1870),
            data_im_out(30) => first_stage_im_out(1934),
            data_im_out(31) => first_stage_im_out(1998)
        );

    ULFFT_PT32_15 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(15),
            data_re_in(1) => data_re_in(79),
            data_re_in(2) => data_re_in(143),
            data_re_in(3) => data_re_in(207),
            data_re_in(4) => data_re_in(271),
            data_re_in(5) => data_re_in(335),
            data_re_in(6) => data_re_in(399),
            data_re_in(7) => data_re_in(463),
            data_re_in(8) => data_re_in(527),
            data_re_in(9) => data_re_in(591),
            data_re_in(10) => data_re_in(655),
            data_re_in(11) => data_re_in(719),
            data_re_in(12) => data_re_in(783),
            data_re_in(13) => data_re_in(847),
            data_re_in(14) => data_re_in(911),
            data_re_in(15) => data_re_in(975),
            data_re_in(16) => data_re_in(1039),
            data_re_in(17) => data_re_in(1103),
            data_re_in(18) => data_re_in(1167),
            data_re_in(19) => data_re_in(1231),
            data_re_in(20) => data_re_in(1295),
            data_re_in(21) => data_re_in(1359),
            data_re_in(22) => data_re_in(1423),
            data_re_in(23) => data_re_in(1487),
            data_re_in(24) => data_re_in(1551),
            data_re_in(25) => data_re_in(1615),
            data_re_in(26) => data_re_in(1679),
            data_re_in(27) => data_re_in(1743),
            data_re_in(28) => data_re_in(1807),
            data_re_in(29) => data_re_in(1871),
            data_re_in(30) => data_re_in(1935),
            data_re_in(31) => data_re_in(1999),
            data_im_in(0) => data_im_in(15),
            data_im_in(1) => data_im_in(79),
            data_im_in(2) => data_im_in(143),
            data_im_in(3) => data_im_in(207),
            data_im_in(4) => data_im_in(271),
            data_im_in(5) => data_im_in(335),
            data_im_in(6) => data_im_in(399),
            data_im_in(7) => data_im_in(463),
            data_im_in(8) => data_im_in(527),
            data_im_in(9) => data_im_in(591),
            data_im_in(10) => data_im_in(655),
            data_im_in(11) => data_im_in(719),
            data_im_in(12) => data_im_in(783),
            data_im_in(13) => data_im_in(847),
            data_im_in(14) => data_im_in(911),
            data_im_in(15) => data_im_in(975),
            data_im_in(16) => data_im_in(1039),
            data_im_in(17) => data_im_in(1103),
            data_im_in(18) => data_im_in(1167),
            data_im_in(19) => data_im_in(1231),
            data_im_in(20) => data_im_in(1295),
            data_im_in(21) => data_im_in(1359),
            data_im_in(22) => data_im_in(1423),
            data_im_in(23) => data_im_in(1487),
            data_im_in(24) => data_im_in(1551),
            data_im_in(25) => data_im_in(1615),
            data_im_in(26) => data_im_in(1679),
            data_im_in(27) => data_im_in(1743),
            data_im_in(28) => data_im_in(1807),
            data_im_in(29) => data_im_in(1871),
            data_im_in(30) => data_im_in(1935),
            data_im_in(31) => data_im_in(1999),
            data_re_out(0) => first_stage_re_out(15),
            data_re_out(1) => first_stage_re_out(79),
            data_re_out(2) => first_stage_re_out(143),
            data_re_out(3) => first_stage_re_out(207),
            data_re_out(4) => first_stage_re_out(271),
            data_re_out(5) => first_stage_re_out(335),
            data_re_out(6) => first_stage_re_out(399),
            data_re_out(7) => first_stage_re_out(463),
            data_re_out(8) => first_stage_re_out(527),
            data_re_out(9) => first_stage_re_out(591),
            data_re_out(10) => first_stage_re_out(655),
            data_re_out(11) => first_stage_re_out(719),
            data_re_out(12) => first_stage_re_out(783),
            data_re_out(13) => first_stage_re_out(847),
            data_re_out(14) => first_stage_re_out(911),
            data_re_out(15) => first_stage_re_out(975),
            data_re_out(16) => first_stage_re_out(1039),
            data_re_out(17) => first_stage_re_out(1103),
            data_re_out(18) => first_stage_re_out(1167),
            data_re_out(19) => first_stage_re_out(1231),
            data_re_out(20) => first_stage_re_out(1295),
            data_re_out(21) => first_stage_re_out(1359),
            data_re_out(22) => first_stage_re_out(1423),
            data_re_out(23) => first_stage_re_out(1487),
            data_re_out(24) => first_stage_re_out(1551),
            data_re_out(25) => first_stage_re_out(1615),
            data_re_out(26) => first_stage_re_out(1679),
            data_re_out(27) => first_stage_re_out(1743),
            data_re_out(28) => first_stage_re_out(1807),
            data_re_out(29) => first_stage_re_out(1871),
            data_re_out(30) => first_stage_re_out(1935),
            data_re_out(31) => first_stage_re_out(1999),
            data_im_out(0) => first_stage_im_out(15),
            data_im_out(1) => first_stage_im_out(79),
            data_im_out(2) => first_stage_im_out(143),
            data_im_out(3) => first_stage_im_out(207),
            data_im_out(4) => first_stage_im_out(271),
            data_im_out(5) => first_stage_im_out(335),
            data_im_out(6) => first_stage_im_out(399),
            data_im_out(7) => first_stage_im_out(463),
            data_im_out(8) => first_stage_im_out(527),
            data_im_out(9) => first_stage_im_out(591),
            data_im_out(10) => first_stage_im_out(655),
            data_im_out(11) => first_stage_im_out(719),
            data_im_out(12) => first_stage_im_out(783),
            data_im_out(13) => first_stage_im_out(847),
            data_im_out(14) => first_stage_im_out(911),
            data_im_out(15) => first_stage_im_out(975),
            data_im_out(16) => first_stage_im_out(1039),
            data_im_out(17) => first_stage_im_out(1103),
            data_im_out(18) => first_stage_im_out(1167),
            data_im_out(19) => first_stage_im_out(1231),
            data_im_out(20) => first_stage_im_out(1295),
            data_im_out(21) => first_stage_im_out(1359),
            data_im_out(22) => first_stage_im_out(1423),
            data_im_out(23) => first_stage_im_out(1487),
            data_im_out(24) => first_stage_im_out(1551),
            data_im_out(25) => first_stage_im_out(1615),
            data_im_out(26) => first_stage_im_out(1679),
            data_im_out(27) => first_stage_im_out(1743),
            data_im_out(28) => first_stage_im_out(1807),
            data_im_out(29) => first_stage_im_out(1871),
            data_im_out(30) => first_stage_im_out(1935),
            data_im_out(31) => first_stage_im_out(1999)
        );

    ULFFT_PT32_16 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(16),
            data_re_in(1) => data_re_in(80),
            data_re_in(2) => data_re_in(144),
            data_re_in(3) => data_re_in(208),
            data_re_in(4) => data_re_in(272),
            data_re_in(5) => data_re_in(336),
            data_re_in(6) => data_re_in(400),
            data_re_in(7) => data_re_in(464),
            data_re_in(8) => data_re_in(528),
            data_re_in(9) => data_re_in(592),
            data_re_in(10) => data_re_in(656),
            data_re_in(11) => data_re_in(720),
            data_re_in(12) => data_re_in(784),
            data_re_in(13) => data_re_in(848),
            data_re_in(14) => data_re_in(912),
            data_re_in(15) => data_re_in(976),
            data_re_in(16) => data_re_in(1040),
            data_re_in(17) => data_re_in(1104),
            data_re_in(18) => data_re_in(1168),
            data_re_in(19) => data_re_in(1232),
            data_re_in(20) => data_re_in(1296),
            data_re_in(21) => data_re_in(1360),
            data_re_in(22) => data_re_in(1424),
            data_re_in(23) => data_re_in(1488),
            data_re_in(24) => data_re_in(1552),
            data_re_in(25) => data_re_in(1616),
            data_re_in(26) => data_re_in(1680),
            data_re_in(27) => data_re_in(1744),
            data_re_in(28) => data_re_in(1808),
            data_re_in(29) => data_re_in(1872),
            data_re_in(30) => data_re_in(1936),
            data_re_in(31) => data_re_in(2000),
            data_im_in(0) => data_im_in(16),
            data_im_in(1) => data_im_in(80),
            data_im_in(2) => data_im_in(144),
            data_im_in(3) => data_im_in(208),
            data_im_in(4) => data_im_in(272),
            data_im_in(5) => data_im_in(336),
            data_im_in(6) => data_im_in(400),
            data_im_in(7) => data_im_in(464),
            data_im_in(8) => data_im_in(528),
            data_im_in(9) => data_im_in(592),
            data_im_in(10) => data_im_in(656),
            data_im_in(11) => data_im_in(720),
            data_im_in(12) => data_im_in(784),
            data_im_in(13) => data_im_in(848),
            data_im_in(14) => data_im_in(912),
            data_im_in(15) => data_im_in(976),
            data_im_in(16) => data_im_in(1040),
            data_im_in(17) => data_im_in(1104),
            data_im_in(18) => data_im_in(1168),
            data_im_in(19) => data_im_in(1232),
            data_im_in(20) => data_im_in(1296),
            data_im_in(21) => data_im_in(1360),
            data_im_in(22) => data_im_in(1424),
            data_im_in(23) => data_im_in(1488),
            data_im_in(24) => data_im_in(1552),
            data_im_in(25) => data_im_in(1616),
            data_im_in(26) => data_im_in(1680),
            data_im_in(27) => data_im_in(1744),
            data_im_in(28) => data_im_in(1808),
            data_im_in(29) => data_im_in(1872),
            data_im_in(30) => data_im_in(1936),
            data_im_in(31) => data_im_in(2000),
            data_re_out(0) => first_stage_re_out(16),
            data_re_out(1) => first_stage_re_out(80),
            data_re_out(2) => first_stage_re_out(144),
            data_re_out(3) => first_stage_re_out(208),
            data_re_out(4) => first_stage_re_out(272),
            data_re_out(5) => first_stage_re_out(336),
            data_re_out(6) => first_stage_re_out(400),
            data_re_out(7) => first_stage_re_out(464),
            data_re_out(8) => first_stage_re_out(528),
            data_re_out(9) => first_stage_re_out(592),
            data_re_out(10) => first_stage_re_out(656),
            data_re_out(11) => first_stage_re_out(720),
            data_re_out(12) => first_stage_re_out(784),
            data_re_out(13) => first_stage_re_out(848),
            data_re_out(14) => first_stage_re_out(912),
            data_re_out(15) => first_stage_re_out(976),
            data_re_out(16) => first_stage_re_out(1040),
            data_re_out(17) => first_stage_re_out(1104),
            data_re_out(18) => first_stage_re_out(1168),
            data_re_out(19) => first_stage_re_out(1232),
            data_re_out(20) => first_stage_re_out(1296),
            data_re_out(21) => first_stage_re_out(1360),
            data_re_out(22) => first_stage_re_out(1424),
            data_re_out(23) => first_stage_re_out(1488),
            data_re_out(24) => first_stage_re_out(1552),
            data_re_out(25) => first_stage_re_out(1616),
            data_re_out(26) => first_stage_re_out(1680),
            data_re_out(27) => first_stage_re_out(1744),
            data_re_out(28) => first_stage_re_out(1808),
            data_re_out(29) => first_stage_re_out(1872),
            data_re_out(30) => first_stage_re_out(1936),
            data_re_out(31) => first_stage_re_out(2000),
            data_im_out(0) => first_stage_im_out(16),
            data_im_out(1) => first_stage_im_out(80),
            data_im_out(2) => first_stage_im_out(144),
            data_im_out(3) => first_stage_im_out(208),
            data_im_out(4) => first_stage_im_out(272),
            data_im_out(5) => first_stage_im_out(336),
            data_im_out(6) => first_stage_im_out(400),
            data_im_out(7) => first_stage_im_out(464),
            data_im_out(8) => first_stage_im_out(528),
            data_im_out(9) => first_stage_im_out(592),
            data_im_out(10) => first_stage_im_out(656),
            data_im_out(11) => first_stage_im_out(720),
            data_im_out(12) => first_stage_im_out(784),
            data_im_out(13) => first_stage_im_out(848),
            data_im_out(14) => first_stage_im_out(912),
            data_im_out(15) => first_stage_im_out(976),
            data_im_out(16) => first_stage_im_out(1040),
            data_im_out(17) => first_stage_im_out(1104),
            data_im_out(18) => first_stage_im_out(1168),
            data_im_out(19) => first_stage_im_out(1232),
            data_im_out(20) => first_stage_im_out(1296),
            data_im_out(21) => first_stage_im_out(1360),
            data_im_out(22) => first_stage_im_out(1424),
            data_im_out(23) => first_stage_im_out(1488),
            data_im_out(24) => first_stage_im_out(1552),
            data_im_out(25) => first_stage_im_out(1616),
            data_im_out(26) => first_stage_im_out(1680),
            data_im_out(27) => first_stage_im_out(1744),
            data_im_out(28) => first_stage_im_out(1808),
            data_im_out(29) => first_stage_im_out(1872),
            data_im_out(30) => first_stage_im_out(1936),
            data_im_out(31) => first_stage_im_out(2000)
        );

    ULFFT_PT32_17 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(17),
            data_re_in(1) => data_re_in(81),
            data_re_in(2) => data_re_in(145),
            data_re_in(3) => data_re_in(209),
            data_re_in(4) => data_re_in(273),
            data_re_in(5) => data_re_in(337),
            data_re_in(6) => data_re_in(401),
            data_re_in(7) => data_re_in(465),
            data_re_in(8) => data_re_in(529),
            data_re_in(9) => data_re_in(593),
            data_re_in(10) => data_re_in(657),
            data_re_in(11) => data_re_in(721),
            data_re_in(12) => data_re_in(785),
            data_re_in(13) => data_re_in(849),
            data_re_in(14) => data_re_in(913),
            data_re_in(15) => data_re_in(977),
            data_re_in(16) => data_re_in(1041),
            data_re_in(17) => data_re_in(1105),
            data_re_in(18) => data_re_in(1169),
            data_re_in(19) => data_re_in(1233),
            data_re_in(20) => data_re_in(1297),
            data_re_in(21) => data_re_in(1361),
            data_re_in(22) => data_re_in(1425),
            data_re_in(23) => data_re_in(1489),
            data_re_in(24) => data_re_in(1553),
            data_re_in(25) => data_re_in(1617),
            data_re_in(26) => data_re_in(1681),
            data_re_in(27) => data_re_in(1745),
            data_re_in(28) => data_re_in(1809),
            data_re_in(29) => data_re_in(1873),
            data_re_in(30) => data_re_in(1937),
            data_re_in(31) => data_re_in(2001),
            data_im_in(0) => data_im_in(17),
            data_im_in(1) => data_im_in(81),
            data_im_in(2) => data_im_in(145),
            data_im_in(3) => data_im_in(209),
            data_im_in(4) => data_im_in(273),
            data_im_in(5) => data_im_in(337),
            data_im_in(6) => data_im_in(401),
            data_im_in(7) => data_im_in(465),
            data_im_in(8) => data_im_in(529),
            data_im_in(9) => data_im_in(593),
            data_im_in(10) => data_im_in(657),
            data_im_in(11) => data_im_in(721),
            data_im_in(12) => data_im_in(785),
            data_im_in(13) => data_im_in(849),
            data_im_in(14) => data_im_in(913),
            data_im_in(15) => data_im_in(977),
            data_im_in(16) => data_im_in(1041),
            data_im_in(17) => data_im_in(1105),
            data_im_in(18) => data_im_in(1169),
            data_im_in(19) => data_im_in(1233),
            data_im_in(20) => data_im_in(1297),
            data_im_in(21) => data_im_in(1361),
            data_im_in(22) => data_im_in(1425),
            data_im_in(23) => data_im_in(1489),
            data_im_in(24) => data_im_in(1553),
            data_im_in(25) => data_im_in(1617),
            data_im_in(26) => data_im_in(1681),
            data_im_in(27) => data_im_in(1745),
            data_im_in(28) => data_im_in(1809),
            data_im_in(29) => data_im_in(1873),
            data_im_in(30) => data_im_in(1937),
            data_im_in(31) => data_im_in(2001),
            data_re_out(0) => first_stage_re_out(17),
            data_re_out(1) => first_stage_re_out(81),
            data_re_out(2) => first_stage_re_out(145),
            data_re_out(3) => first_stage_re_out(209),
            data_re_out(4) => first_stage_re_out(273),
            data_re_out(5) => first_stage_re_out(337),
            data_re_out(6) => first_stage_re_out(401),
            data_re_out(7) => first_stage_re_out(465),
            data_re_out(8) => first_stage_re_out(529),
            data_re_out(9) => first_stage_re_out(593),
            data_re_out(10) => first_stage_re_out(657),
            data_re_out(11) => first_stage_re_out(721),
            data_re_out(12) => first_stage_re_out(785),
            data_re_out(13) => first_stage_re_out(849),
            data_re_out(14) => first_stage_re_out(913),
            data_re_out(15) => first_stage_re_out(977),
            data_re_out(16) => first_stage_re_out(1041),
            data_re_out(17) => first_stage_re_out(1105),
            data_re_out(18) => first_stage_re_out(1169),
            data_re_out(19) => first_stage_re_out(1233),
            data_re_out(20) => first_stage_re_out(1297),
            data_re_out(21) => first_stage_re_out(1361),
            data_re_out(22) => first_stage_re_out(1425),
            data_re_out(23) => first_stage_re_out(1489),
            data_re_out(24) => first_stage_re_out(1553),
            data_re_out(25) => first_stage_re_out(1617),
            data_re_out(26) => first_stage_re_out(1681),
            data_re_out(27) => first_stage_re_out(1745),
            data_re_out(28) => first_stage_re_out(1809),
            data_re_out(29) => first_stage_re_out(1873),
            data_re_out(30) => first_stage_re_out(1937),
            data_re_out(31) => first_stage_re_out(2001),
            data_im_out(0) => first_stage_im_out(17),
            data_im_out(1) => first_stage_im_out(81),
            data_im_out(2) => first_stage_im_out(145),
            data_im_out(3) => first_stage_im_out(209),
            data_im_out(4) => first_stage_im_out(273),
            data_im_out(5) => first_stage_im_out(337),
            data_im_out(6) => first_stage_im_out(401),
            data_im_out(7) => first_stage_im_out(465),
            data_im_out(8) => first_stage_im_out(529),
            data_im_out(9) => first_stage_im_out(593),
            data_im_out(10) => first_stage_im_out(657),
            data_im_out(11) => first_stage_im_out(721),
            data_im_out(12) => first_stage_im_out(785),
            data_im_out(13) => first_stage_im_out(849),
            data_im_out(14) => first_stage_im_out(913),
            data_im_out(15) => first_stage_im_out(977),
            data_im_out(16) => first_stage_im_out(1041),
            data_im_out(17) => first_stage_im_out(1105),
            data_im_out(18) => first_stage_im_out(1169),
            data_im_out(19) => first_stage_im_out(1233),
            data_im_out(20) => first_stage_im_out(1297),
            data_im_out(21) => first_stage_im_out(1361),
            data_im_out(22) => first_stage_im_out(1425),
            data_im_out(23) => first_stage_im_out(1489),
            data_im_out(24) => first_stage_im_out(1553),
            data_im_out(25) => first_stage_im_out(1617),
            data_im_out(26) => first_stage_im_out(1681),
            data_im_out(27) => first_stage_im_out(1745),
            data_im_out(28) => first_stage_im_out(1809),
            data_im_out(29) => first_stage_im_out(1873),
            data_im_out(30) => first_stage_im_out(1937),
            data_im_out(31) => first_stage_im_out(2001)
        );

    ULFFT_PT32_18 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(18),
            data_re_in(1) => data_re_in(82),
            data_re_in(2) => data_re_in(146),
            data_re_in(3) => data_re_in(210),
            data_re_in(4) => data_re_in(274),
            data_re_in(5) => data_re_in(338),
            data_re_in(6) => data_re_in(402),
            data_re_in(7) => data_re_in(466),
            data_re_in(8) => data_re_in(530),
            data_re_in(9) => data_re_in(594),
            data_re_in(10) => data_re_in(658),
            data_re_in(11) => data_re_in(722),
            data_re_in(12) => data_re_in(786),
            data_re_in(13) => data_re_in(850),
            data_re_in(14) => data_re_in(914),
            data_re_in(15) => data_re_in(978),
            data_re_in(16) => data_re_in(1042),
            data_re_in(17) => data_re_in(1106),
            data_re_in(18) => data_re_in(1170),
            data_re_in(19) => data_re_in(1234),
            data_re_in(20) => data_re_in(1298),
            data_re_in(21) => data_re_in(1362),
            data_re_in(22) => data_re_in(1426),
            data_re_in(23) => data_re_in(1490),
            data_re_in(24) => data_re_in(1554),
            data_re_in(25) => data_re_in(1618),
            data_re_in(26) => data_re_in(1682),
            data_re_in(27) => data_re_in(1746),
            data_re_in(28) => data_re_in(1810),
            data_re_in(29) => data_re_in(1874),
            data_re_in(30) => data_re_in(1938),
            data_re_in(31) => data_re_in(2002),
            data_im_in(0) => data_im_in(18),
            data_im_in(1) => data_im_in(82),
            data_im_in(2) => data_im_in(146),
            data_im_in(3) => data_im_in(210),
            data_im_in(4) => data_im_in(274),
            data_im_in(5) => data_im_in(338),
            data_im_in(6) => data_im_in(402),
            data_im_in(7) => data_im_in(466),
            data_im_in(8) => data_im_in(530),
            data_im_in(9) => data_im_in(594),
            data_im_in(10) => data_im_in(658),
            data_im_in(11) => data_im_in(722),
            data_im_in(12) => data_im_in(786),
            data_im_in(13) => data_im_in(850),
            data_im_in(14) => data_im_in(914),
            data_im_in(15) => data_im_in(978),
            data_im_in(16) => data_im_in(1042),
            data_im_in(17) => data_im_in(1106),
            data_im_in(18) => data_im_in(1170),
            data_im_in(19) => data_im_in(1234),
            data_im_in(20) => data_im_in(1298),
            data_im_in(21) => data_im_in(1362),
            data_im_in(22) => data_im_in(1426),
            data_im_in(23) => data_im_in(1490),
            data_im_in(24) => data_im_in(1554),
            data_im_in(25) => data_im_in(1618),
            data_im_in(26) => data_im_in(1682),
            data_im_in(27) => data_im_in(1746),
            data_im_in(28) => data_im_in(1810),
            data_im_in(29) => data_im_in(1874),
            data_im_in(30) => data_im_in(1938),
            data_im_in(31) => data_im_in(2002),
            data_re_out(0) => first_stage_re_out(18),
            data_re_out(1) => first_stage_re_out(82),
            data_re_out(2) => first_stage_re_out(146),
            data_re_out(3) => first_stage_re_out(210),
            data_re_out(4) => first_stage_re_out(274),
            data_re_out(5) => first_stage_re_out(338),
            data_re_out(6) => first_stage_re_out(402),
            data_re_out(7) => first_stage_re_out(466),
            data_re_out(8) => first_stage_re_out(530),
            data_re_out(9) => first_stage_re_out(594),
            data_re_out(10) => first_stage_re_out(658),
            data_re_out(11) => first_stage_re_out(722),
            data_re_out(12) => first_stage_re_out(786),
            data_re_out(13) => first_stage_re_out(850),
            data_re_out(14) => first_stage_re_out(914),
            data_re_out(15) => first_stage_re_out(978),
            data_re_out(16) => first_stage_re_out(1042),
            data_re_out(17) => first_stage_re_out(1106),
            data_re_out(18) => first_stage_re_out(1170),
            data_re_out(19) => first_stage_re_out(1234),
            data_re_out(20) => first_stage_re_out(1298),
            data_re_out(21) => first_stage_re_out(1362),
            data_re_out(22) => first_stage_re_out(1426),
            data_re_out(23) => first_stage_re_out(1490),
            data_re_out(24) => first_stage_re_out(1554),
            data_re_out(25) => first_stage_re_out(1618),
            data_re_out(26) => first_stage_re_out(1682),
            data_re_out(27) => first_stage_re_out(1746),
            data_re_out(28) => first_stage_re_out(1810),
            data_re_out(29) => first_stage_re_out(1874),
            data_re_out(30) => first_stage_re_out(1938),
            data_re_out(31) => first_stage_re_out(2002),
            data_im_out(0) => first_stage_im_out(18),
            data_im_out(1) => first_stage_im_out(82),
            data_im_out(2) => first_stage_im_out(146),
            data_im_out(3) => first_stage_im_out(210),
            data_im_out(4) => first_stage_im_out(274),
            data_im_out(5) => first_stage_im_out(338),
            data_im_out(6) => first_stage_im_out(402),
            data_im_out(7) => first_stage_im_out(466),
            data_im_out(8) => first_stage_im_out(530),
            data_im_out(9) => first_stage_im_out(594),
            data_im_out(10) => first_stage_im_out(658),
            data_im_out(11) => first_stage_im_out(722),
            data_im_out(12) => first_stage_im_out(786),
            data_im_out(13) => first_stage_im_out(850),
            data_im_out(14) => first_stage_im_out(914),
            data_im_out(15) => first_stage_im_out(978),
            data_im_out(16) => first_stage_im_out(1042),
            data_im_out(17) => first_stage_im_out(1106),
            data_im_out(18) => first_stage_im_out(1170),
            data_im_out(19) => first_stage_im_out(1234),
            data_im_out(20) => first_stage_im_out(1298),
            data_im_out(21) => first_stage_im_out(1362),
            data_im_out(22) => first_stage_im_out(1426),
            data_im_out(23) => first_stage_im_out(1490),
            data_im_out(24) => first_stage_im_out(1554),
            data_im_out(25) => first_stage_im_out(1618),
            data_im_out(26) => first_stage_im_out(1682),
            data_im_out(27) => first_stage_im_out(1746),
            data_im_out(28) => first_stage_im_out(1810),
            data_im_out(29) => first_stage_im_out(1874),
            data_im_out(30) => first_stage_im_out(1938),
            data_im_out(31) => first_stage_im_out(2002)
        );

    ULFFT_PT32_19 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(19),
            data_re_in(1) => data_re_in(83),
            data_re_in(2) => data_re_in(147),
            data_re_in(3) => data_re_in(211),
            data_re_in(4) => data_re_in(275),
            data_re_in(5) => data_re_in(339),
            data_re_in(6) => data_re_in(403),
            data_re_in(7) => data_re_in(467),
            data_re_in(8) => data_re_in(531),
            data_re_in(9) => data_re_in(595),
            data_re_in(10) => data_re_in(659),
            data_re_in(11) => data_re_in(723),
            data_re_in(12) => data_re_in(787),
            data_re_in(13) => data_re_in(851),
            data_re_in(14) => data_re_in(915),
            data_re_in(15) => data_re_in(979),
            data_re_in(16) => data_re_in(1043),
            data_re_in(17) => data_re_in(1107),
            data_re_in(18) => data_re_in(1171),
            data_re_in(19) => data_re_in(1235),
            data_re_in(20) => data_re_in(1299),
            data_re_in(21) => data_re_in(1363),
            data_re_in(22) => data_re_in(1427),
            data_re_in(23) => data_re_in(1491),
            data_re_in(24) => data_re_in(1555),
            data_re_in(25) => data_re_in(1619),
            data_re_in(26) => data_re_in(1683),
            data_re_in(27) => data_re_in(1747),
            data_re_in(28) => data_re_in(1811),
            data_re_in(29) => data_re_in(1875),
            data_re_in(30) => data_re_in(1939),
            data_re_in(31) => data_re_in(2003),
            data_im_in(0) => data_im_in(19),
            data_im_in(1) => data_im_in(83),
            data_im_in(2) => data_im_in(147),
            data_im_in(3) => data_im_in(211),
            data_im_in(4) => data_im_in(275),
            data_im_in(5) => data_im_in(339),
            data_im_in(6) => data_im_in(403),
            data_im_in(7) => data_im_in(467),
            data_im_in(8) => data_im_in(531),
            data_im_in(9) => data_im_in(595),
            data_im_in(10) => data_im_in(659),
            data_im_in(11) => data_im_in(723),
            data_im_in(12) => data_im_in(787),
            data_im_in(13) => data_im_in(851),
            data_im_in(14) => data_im_in(915),
            data_im_in(15) => data_im_in(979),
            data_im_in(16) => data_im_in(1043),
            data_im_in(17) => data_im_in(1107),
            data_im_in(18) => data_im_in(1171),
            data_im_in(19) => data_im_in(1235),
            data_im_in(20) => data_im_in(1299),
            data_im_in(21) => data_im_in(1363),
            data_im_in(22) => data_im_in(1427),
            data_im_in(23) => data_im_in(1491),
            data_im_in(24) => data_im_in(1555),
            data_im_in(25) => data_im_in(1619),
            data_im_in(26) => data_im_in(1683),
            data_im_in(27) => data_im_in(1747),
            data_im_in(28) => data_im_in(1811),
            data_im_in(29) => data_im_in(1875),
            data_im_in(30) => data_im_in(1939),
            data_im_in(31) => data_im_in(2003),
            data_re_out(0) => first_stage_re_out(19),
            data_re_out(1) => first_stage_re_out(83),
            data_re_out(2) => first_stage_re_out(147),
            data_re_out(3) => first_stage_re_out(211),
            data_re_out(4) => first_stage_re_out(275),
            data_re_out(5) => first_stage_re_out(339),
            data_re_out(6) => first_stage_re_out(403),
            data_re_out(7) => first_stage_re_out(467),
            data_re_out(8) => first_stage_re_out(531),
            data_re_out(9) => first_stage_re_out(595),
            data_re_out(10) => first_stage_re_out(659),
            data_re_out(11) => first_stage_re_out(723),
            data_re_out(12) => first_stage_re_out(787),
            data_re_out(13) => first_stage_re_out(851),
            data_re_out(14) => first_stage_re_out(915),
            data_re_out(15) => first_stage_re_out(979),
            data_re_out(16) => first_stage_re_out(1043),
            data_re_out(17) => first_stage_re_out(1107),
            data_re_out(18) => first_stage_re_out(1171),
            data_re_out(19) => first_stage_re_out(1235),
            data_re_out(20) => first_stage_re_out(1299),
            data_re_out(21) => first_stage_re_out(1363),
            data_re_out(22) => first_stage_re_out(1427),
            data_re_out(23) => first_stage_re_out(1491),
            data_re_out(24) => first_stage_re_out(1555),
            data_re_out(25) => first_stage_re_out(1619),
            data_re_out(26) => first_stage_re_out(1683),
            data_re_out(27) => first_stage_re_out(1747),
            data_re_out(28) => first_stage_re_out(1811),
            data_re_out(29) => first_stage_re_out(1875),
            data_re_out(30) => first_stage_re_out(1939),
            data_re_out(31) => first_stage_re_out(2003),
            data_im_out(0) => first_stage_im_out(19),
            data_im_out(1) => first_stage_im_out(83),
            data_im_out(2) => first_stage_im_out(147),
            data_im_out(3) => first_stage_im_out(211),
            data_im_out(4) => first_stage_im_out(275),
            data_im_out(5) => first_stage_im_out(339),
            data_im_out(6) => first_stage_im_out(403),
            data_im_out(7) => first_stage_im_out(467),
            data_im_out(8) => first_stage_im_out(531),
            data_im_out(9) => first_stage_im_out(595),
            data_im_out(10) => first_stage_im_out(659),
            data_im_out(11) => first_stage_im_out(723),
            data_im_out(12) => first_stage_im_out(787),
            data_im_out(13) => first_stage_im_out(851),
            data_im_out(14) => first_stage_im_out(915),
            data_im_out(15) => first_stage_im_out(979),
            data_im_out(16) => first_stage_im_out(1043),
            data_im_out(17) => first_stage_im_out(1107),
            data_im_out(18) => first_stage_im_out(1171),
            data_im_out(19) => first_stage_im_out(1235),
            data_im_out(20) => first_stage_im_out(1299),
            data_im_out(21) => first_stage_im_out(1363),
            data_im_out(22) => first_stage_im_out(1427),
            data_im_out(23) => first_stage_im_out(1491),
            data_im_out(24) => first_stage_im_out(1555),
            data_im_out(25) => first_stage_im_out(1619),
            data_im_out(26) => first_stage_im_out(1683),
            data_im_out(27) => first_stage_im_out(1747),
            data_im_out(28) => first_stage_im_out(1811),
            data_im_out(29) => first_stage_im_out(1875),
            data_im_out(30) => first_stage_im_out(1939),
            data_im_out(31) => first_stage_im_out(2003)
        );

    ULFFT_PT32_20 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(20),
            data_re_in(1) => data_re_in(84),
            data_re_in(2) => data_re_in(148),
            data_re_in(3) => data_re_in(212),
            data_re_in(4) => data_re_in(276),
            data_re_in(5) => data_re_in(340),
            data_re_in(6) => data_re_in(404),
            data_re_in(7) => data_re_in(468),
            data_re_in(8) => data_re_in(532),
            data_re_in(9) => data_re_in(596),
            data_re_in(10) => data_re_in(660),
            data_re_in(11) => data_re_in(724),
            data_re_in(12) => data_re_in(788),
            data_re_in(13) => data_re_in(852),
            data_re_in(14) => data_re_in(916),
            data_re_in(15) => data_re_in(980),
            data_re_in(16) => data_re_in(1044),
            data_re_in(17) => data_re_in(1108),
            data_re_in(18) => data_re_in(1172),
            data_re_in(19) => data_re_in(1236),
            data_re_in(20) => data_re_in(1300),
            data_re_in(21) => data_re_in(1364),
            data_re_in(22) => data_re_in(1428),
            data_re_in(23) => data_re_in(1492),
            data_re_in(24) => data_re_in(1556),
            data_re_in(25) => data_re_in(1620),
            data_re_in(26) => data_re_in(1684),
            data_re_in(27) => data_re_in(1748),
            data_re_in(28) => data_re_in(1812),
            data_re_in(29) => data_re_in(1876),
            data_re_in(30) => data_re_in(1940),
            data_re_in(31) => data_re_in(2004),
            data_im_in(0) => data_im_in(20),
            data_im_in(1) => data_im_in(84),
            data_im_in(2) => data_im_in(148),
            data_im_in(3) => data_im_in(212),
            data_im_in(4) => data_im_in(276),
            data_im_in(5) => data_im_in(340),
            data_im_in(6) => data_im_in(404),
            data_im_in(7) => data_im_in(468),
            data_im_in(8) => data_im_in(532),
            data_im_in(9) => data_im_in(596),
            data_im_in(10) => data_im_in(660),
            data_im_in(11) => data_im_in(724),
            data_im_in(12) => data_im_in(788),
            data_im_in(13) => data_im_in(852),
            data_im_in(14) => data_im_in(916),
            data_im_in(15) => data_im_in(980),
            data_im_in(16) => data_im_in(1044),
            data_im_in(17) => data_im_in(1108),
            data_im_in(18) => data_im_in(1172),
            data_im_in(19) => data_im_in(1236),
            data_im_in(20) => data_im_in(1300),
            data_im_in(21) => data_im_in(1364),
            data_im_in(22) => data_im_in(1428),
            data_im_in(23) => data_im_in(1492),
            data_im_in(24) => data_im_in(1556),
            data_im_in(25) => data_im_in(1620),
            data_im_in(26) => data_im_in(1684),
            data_im_in(27) => data_im_in(1748),
            data_im_in(28) => data_im_in(1812),
            data_im_in(29) => data_im_in(1876),
            data_im_in(30) => data_im_in(1940),
            data_im_in(31) => data_im_in(2004),
            data_re_out(0) => first_stage_re_out(20),
            data_re_out(1) => first_stage_re_out(84),
            data_re_out(2) => first_stage_re_out(148),
            data_re_out(3) => first_stage_re_out(212),
            data_re_out(4) => first_stage_re_out(276),
            data_re_out(5) => first_stage_re_out(340),
            data_re_out(6) => first_stage_re_out(404),
            data_re_out(7) => first_stage_re_out(468),
            data_re_out(8) => first_stage_re_out(532),
            data_re_out(9) => first_stage_re_out(596),
            data_re_out(10) => first_stage_re_out(660),
            data_re_out(11) => first_stage_re_out(724),
            data_re_out(12) => first_stage_re_out(788),
            data_re_out(13) => first_stage_re_out(852),
            data_re_out(14) => first_stage_re_out(916),
            data_re_out(15) => first_stage_re_out(980),
            data_re_out(16) => first_stage_re_out(1044),
            data_re_out(17) => first_stage_re_out(1108),
            data_re_out(18) => first_stage_re_out(1172),
            data_re_out(19) => first_stage_re_out(1236),
            data_re_out(20) => first_stage_re_out(1300),
            data_re_out(21) => first_stage_re_out(1364),
            data_re_out(22) => first_stage_re_out(1428),
            data_re_out(23) => first_stage_re_out(1492),
            data_re_out(24) => first_stage_re_out(1556),
            data_re_out(25) => first_stage_re_out(1620),
            data_re_out(26) => first_stage_re_out(1684),
            data_re_out(27) => first_stage_re_out(1748),
            data_re_out(28) => first_stage_re_out(1812),
            data_re_out(29) => first_stage_re_out(1876),
            data_re_out(30) => first_stage_re_out(1940),
            data_re_out(31) => first_stage_re_out(2004),
            data_im_out(0) => first_stage_im_out(20),
            data_im_out(1) => first_stage_im_out(84),
            data_im_out(2) => first_stage_im_out(148),
            data_im_out(3) => first_stage_im_out(212),
            data_im_out(4) => first_stage_im_out(276),
            data_im_out(5) => first_stage_im_out(340),
            data_im_out(6) => first_stage_im_out(404),
            data_im_out(7) => first_stage_im_out(468),
            data_im_out(8) => first_stage_im_out(532),
            data_im_out(9) => first_stage_im_out(596),
            data_im_out(10) => first_stage_im_out(660),
            data_im_out(11) => first_stage_im_out(724),
            data_im_out(12) => first_stage_im_out(788),
            data_im_out(13) => first_stage_im_out(852),
            data_im_out(14) => first_stage_im_out(916),
            data_im_out(15) => first_stage_im_out(980),
            data_im_out(16) => first_stage_im_out(1044),
            data_im_out(17) => first_stage_im_out(1108),
            data_im_out(18) => first_stage_im_out(1172),
            data_im_out(19) => first_stage_im_out(1236),
            data_im_out(20) => first_stage_im_out(1300),
            data_im_out(21) => first_stage_im_out(1364),
            data_im_out(22) => first_stage_im_out(1428),
            data_im_out(23) => first_stage_im_out(1492),
            data_im_out(24) => first_stage_im_out(1556),
            data_im_out(25) => first_stage_im_out(1620),
            data_im_out(26) => first_stage_im_out(1684),
            data_im_out(27) => first_stage_im_out(1748),
            data_im_out(28) => first_stage_im_out(1812),
            data_im_out(29) => first_stage_im_out(1876),
            data_im_out(30) => first_stage_im_out(1940),
            data_im_out(31) => first_stage_im_out(2004)
        );

    ULFFT_PT32_21 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(21),
            data_re_in(1) => data_re_in(85),
            data_re_in(2) => data_re_in(149),
            data_re_in(3) => data_re_in(213),
            data_re_in(4) => data_re_in(277),
            data_re_in(5) => data_re_in(341),
            data_re_in(6) => data_re_in(405),
            data_re_in(7) => data_re_in(469),
            data_re_in(8) => data_re_in(533),
            data_re_in(9) => data_re_in(597),
            data_re_in(10) => data_re_in(661),
            data_re_in(11) => data_re_in(725),
            data_re_in(12) => data_re_in(789),
            data_re_in(13) => data_re_in(853),
            data_re_in(14) => data_re_in(917),
            data_re_in(15) => data_re_in(981),
            data_re_in(16) => data_re_in(1045),
            data_re_in(17) => data_re_in(1109),
            data_re_in(18) => data_re_in(1173),
            data_re_in(19) => data_re_in(1237),
            data_re_in(20) => data_re_in(1301),
            data_re_in(21) => data_re_in(1365),
            data_re_in(22) => data_re_in(1429),
            data_re_in(23) => data_re_in(1493),
            data_re_in(24) => data_re_in(1557),
            data_re_in(25) => data_re_in(1621),
            data_re_in(26) => data_re_in(1685),
            data_re_in(27) => data_re_in(1749),
            data_re_in(28) => data_re_in(1813),
            data_re_in(29) => data_re_in(1877),
            data_re_in(30) => data_re_in(1941),
            data_re_in(31) => data_re_in(2005),
            data_im_in(0) => data_im_in(21),
            data_im_in(1) => data_im_in(85),
            data_im_in(2) => data_im_in(149),
            data_im_in(3) => data_im_in(213),
            data_im_in(4) => data_im_in(277),
            data_im_in(5) => data_im_in(341),
            data_im_in(6) => data_im_in(405),
            data_im_in(7) => data_im_in(469),
            data_im_in(8) => data_im_in(533),
            data_im_in(9) => data_im_in(597),
            data_im_in(10) => data_im_in(661),
            data_im_in(11) => data_im_in(725),
            data_im_in(12) => data_im_in(789),
            data_im_in(13) => data_im_in(853),
            data_im_in(14) => data_im_in(917),
            data_im_in(15) => data_im_in(981),
            data_im_in(16) => data_im_in(1045),
            data_im_in(17) => data_im_in(1109),
            data_im_in(18) => data_im_in(1173),
            data_im_in(19) => data_im_in(1237),
            data_im_in(20) => data_im_in(1301),
            data_im_in(21) => data_im_in(1365),
            data_im_in(22) => data_im_in(1429),
            data_im_in(23) => data_im_in(1493),
            data_im_in(24) => data_im_in(1557),
            data_im_in(25) => data_im_in(1621),
            data_im_in(26) => data_im_in(1685),
            data_im_in(27) => data_im_in(1749),
            data_im_in(28) => data_im_in(1813),
            data_im_in(29) => data_im_in(1877),
            data_im_in(30) => data_im_in(1941),
            data_im_in(31) => data_im_in(2005),
            data_re_out(0) => first_stage_re_out(21),
            data_re_out(1) => first_stage_re_out(85),
            data_re_out(2) => first_stage_re_out(149),
            data_re_out(3) => first_stage_re_out(213),
            data_re_out(4) => first_stage_re_out(277),
            data_re_out(5) => first_stage_re_out(341),
            data_re_out(6) => first_stage_re_out(405),
            data_re_out(7) => first_stage_re_out(469),
            data_re_out(8) => first_stage_re_out(533),
            data_re_out(9) => first_stage_re_out(597),
            data_re_out(10) => first_stage_re_out(661),
            data_re_out(11) => first_stage_re_out(725),
            data_re_out(12) => first_stage_re_out(789),
            data_re_out(13) => first_stage_re_out(853),
            data_re_out(14) => first_stage_re_out(917),
            data_re_out(15) => first_stage_re_out(981),
            data_re_out(16) => first_stage_re_out(1045),
            data_re_out(17) => first_stage_re_out(1109),
            data_re_out(18) => first_stage_re_out(1173),
            data_re_out(19) => first_stage_re_out(1237),
            data_re_out(20) => first_stage_re_out(1301),
            data_re_out(21) => first_stage_re_out(1365),
            data_re_out(22) => first_stage_re_out(1429),
            data_re_out(23) => first_stage_re_out(1493),
            data_re_out(24) => first_stage_re_out(1557),
            data_re_out(25) => first_stage_re_out(1621),
            data_re_out(26) => first_stage_re_out(1685),
            data_re_out(27) => first_stage_re_out(1749),
            data_re_out(28) => first_stage_re_out(1813),
            data_re_out(29) => first_stage_re_out(1877),
            data_re_out(30) => first_stage_re_out(1941),
            data_re_out(31) => first_stage_re_out(2005),
            data_im_out(0) => first_stage_im_out(21),
            data_im_out(1) => first_stage_im_out(85),
            data_im_out(2) => first_stage_im_out(149),
            data_im_out(3) => first_stage_im_out(213),
            data_im_out(4) => first_stage_im_out(277),
            data_im_out(5) => first_stage_im_out(341),
            data_im_out(6) => first_stage_im_out(405),
            data_im_out(7) => first_stage_im_out(469),
            data_im_out(8) => first_stage_im_out(533),
            data_im_out(9) => first_stage_im_out(597),
            data_im_out(10) => first_stage_im_out(661),
            data_im_out(11) => first_stage_im_out(725),
            data_im_out(12) => first_stage_im_out(789),
            data_im_out(13) => first_stage_im_out(853),
            data_im_out(14) => first_stage_im_out(917),
            data_im_out(15) => first_stage_im_out(981),
            data_im_out(16) => first_stage_im_out(1045),
            data_im_out(17) => first_stage_im_out(1109),
            data_im_out(18) => first_stage_im_out(1173),
            data_im_out(19) => first_stage_im_out(1237),
            data_im_out(20) => first_stage_im_out(1301),
            data_im_out(21) => first_stage_im_out(1365),
            data_im_out(22) => first_stage_im_out(1429),
            data_im_out(23) => first_stage_im_out(1493),
            data_im_out(24) => first_stage_im_out(1557),
            data_im_out(25) => first_stage_im_out(1621),
            data_im_out(26) => first_stage_im_out(1685),
            data_im_out(27) => first_stage_im_out(1749),
            data_im_out(28) => first_stage_im_out(1813),
            data_im_out(29) => first_stage_im_out(1877),
            data_im_out(30) => first_stage_im_out(1941),
            data_im_out(31) => first_stage_im_out(2005)
        );

    ULFFT_PT32_22 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(22),
            data_re_in(1) => data_re_in(86),
            data_re_in(2) => data_re_in(150),
            data_re_in(3) => data_re_in(214),
            data_re_in(4) => data_re_in(278),
            data_re_in(5) => data_re_in(342),
            data_re_in(6) => data_re_in(406),
            data_re_in(7) => data_re_in(470),
            data_re_in(8) => data_re_in(534),
            data_re_in(9) => data_re_in(598),
            data_re_in(10) => data_re_in(662),
            data_re_in(11) => data_re_in(726),
            data_re_in(12) => data_re_in(790),
            data_re_in(13) => data_re_in(854),
            data_re_in(14) => data_re_in(918),
            data_re_in(15) => data_re_in(982),
            data_re_in(16) => data_re_in(1046),
            data_re_in(17) => data_re_in(1110),
            data_re_in(18) => data_re_in(1174),
            data_re_in(19) => data_re_in(1238),
            data_re_in(20) => data_re_in(1302),
            data_re_in(21) => data_re_in(1366),
            data_re_in(22) => data_re_in(1430),
            data_re_in(23) => data_re_in(1494),
            data_re_in(24) => data_re_in(1558),
            data_re_in(25) => data_re_in(1622),
            data_re_in(26) => data_re_in(1686),
            data_re_in(27) => data_re_in(1750),
            data_re_in(28) => data_re_in(1814),
            data_re_in(29) => data_re_in(1878),
            data_re_in(30) => data_re_in(1942),
            data_re_in(31) => data_re_in(2006),
            data_im_in(0) => data_im_in(22),
            data_im_in(1) => data_im_in(86),
            data_im_in(2) => data_im_in(150),
            data_im_in(3) => data_im_in(214),
            data_im_in(4) => data_im_in(278),
            data_im_in(5) => data_im_in(342),
            data_im_in(6) => data_im_in(406),
            data_im_in(7) => data_im_in(470),
            data_im_in(8) => data_im_in(534),
            data_im_in(9) => data_im_in(598),
            data_im_in(10) => data_im_in(662),
            data_im_in(11) => data_im_in(726),
            data_im_in(12) => data_im_in(790),
            data_im_in(13) => data_im_in(854),
            data_im_in(14) => data_im_in(918),
            data_im_in(15) => data_im_in(982),
            data_im_in(16) => data_im_in(1046),
            data_im_in(17) => data_im_in(1110),
            data_im_in(18) => data_im_in(1174),
            data_im_in(19) => data_im_in(1238),
            data_im_in(20) => data_im_in(1302),
            data_im_in(21) => data_im_in(1366),
            data_im_in(22) => data_im_in(1430),
            data_im_in(23) => data_im_in(1494),
            data_im_in(24) => data_im_in(1558),
            data_im_in(25) => data_im_in(1622),
            data_im_in(26) => data_im_in(1686),
            data_im_in(27) => data_im_in(1750),
            data_im_in(28) => data_im_in(1814),
            data_im_in(29) => data_im_in(1878),
            data_im_in(30) => data_im_in(1942),
            data_im_in(31) => data_im_in(2006),
            data_re_out(0) => first_stage_re_out(22),
            data_re_out(1) => first_stage_re_out(86),
            data_re_out(2) => first_stage_re_out(150),
            data_re_out(3) => first_stage_re_out(214),
            data_re_out(4) => first_stage_re_out(278),
            data_re_out(5) => first_stage_re_out(342),
            data_re_out(6) => first_stage_re_out(406),
            data_re_out(7) => first_stage_re_out(470),
            data_re_out(8) => first_stage_re_out(534),
            data_re_out(9) => first_stage_re_out(598),
            data_re_out(10) => first_stage_re_out(662),
            data_re_out(11) => first_stage_re_out(726),
            data_re_out(12) => first_stage_re_out(790),
            data_re_out(13) => first_stage_re_out(854),
            data_re_out(14) => first_stage_re_out(918),
            data_re_out(15) => first_stage_re_out(982),
            data_re_out(16) => first_stage_re_out(1046),
            data_re_out(17) => first_stage_re_out(1110),
            data_re_out(18) => first_stage_re_out(1174),
            data_re_out(19) => first_stage_re_out(1238),
            data_re_out(20) => first_stage_re_out(1302),
            data_re_out(21) => first_stage_re_out(1366),
            data_re_out(22) => first_stage_re_out(1430),
            data_re_out(23) => first_stage_re_out(1494),
            data_re_out(24) => first_stage_re_out(1558),
            data_re_out(25) => first_stage_re_out(1622),
            data_re_out(26) => first_stage_re_out(1686),
            data_re_out(27) => first_stage_re_out(1750),
            data_re_out(28) => first_stage_re_out(1814),
            data_re_out(29) => first_stage_re_out(1878),
            data_re_out(30) => first_stage_re_out(1942),
            data_re_out(31) => first_stage_re_out(2006),
            data_im_out(0) => first_stage_im_out(22),
            data_im_out(1) => first_stage_im_out(86),
            data_im_out(2) => first_stage_im_out(150),
            data_im_out(3) => first_stage_im_out(214),
            data_im_out(4) => first_stage_im_out(278),
            data_im_out(5) => first_stage_im_out(342),
            data_im_out(6) => first_stage_im_out(406),
            data_im_out(7) => first_stage_im_out(470),
            data_im_out(8) => first_stage_im_out(534),
            data_im_out(9) => first_stage_im_out(598),
            data_im_out(10) => first_stage_im_out(662),
            data_im_out(11) => first_stage_im_out(726),
            data_im_out(12) => first_stage_im_out(790),
            data_im_out(13) => first_stage_im_out(854),
            data_im_out(14) => first_stage_im_out(918),
            data_im_out(15) => first_stage_im_out(982),
            data_im_out(16) => first_stage_im_out(1046),
            data_im_out(17) => first_stage_im_out(1110),
            data_im_out(18) => first_stage_im_out(1174),
            data_im_out(19) => first_stage_im_out(1238),
            data_im_out(20) => first_stage_im_out(1302),
            data_im_out(21) => first_stage_im_out(1366),
            data_im_out(22) => first_stage_im_out(1430),
            data_im_out(23) => first_stage_im_out(1494),
            data_im_out(24) => first_stage_im_out(1558),
            data_im_out(25) => first_stage_im_out(1622),
            data_im_out(26) => first_stage_im_out(1686),
            data_im_out(27) => first_stage_im_out(1750),
            data_im_out(28) => first_stage_im_out(1814),
            data_im_out(29) => first_stage_im_out(1878),
            data_im_out(30) => first_stage_im_out(1942),
            data_im_out(31) => first_stage_im_out(2006)
        );

    ULFFT_PT32_23 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(23),
            data_re_in(1) => data_re_in(87),
            data_re_in(2) => data_re_in(151),
            data_re_in(3) => data_re_in(215),
            data_re_in(4) => data_re_in(279),
            data_re_in(5) => data_re_in(343),
            data_re_in(6) => data_re_in(407),
            data_re_in(7) => data_re_in(471),
            data_re_in(8) => data_re_in(535),
            data_re_in(9) => data_re_in(599),
            data_re_in(10) => data_re_in(663),
            data_re_in(11) => data_re_in(727),
            data_re_in(12) => data_re_in(791),
            data_re_in(13) => data_re_in(855),
            data_re_in(14) => data_re_in(919),
            data_re_in(15) => data_re_in(983),
            data_re_in(16) => data_re_in(1047),
            data_re_in(17) => data_re_in(1111),
            data_re_in(18) => data_re_in(1175),
            data_re_in(19) => data_re_in(1239),
            data_re_in(20) => data_re_in(1303),
            data_re_in(21) => data_re_in(1367),
            data_re_in(22) => data_re_in(1431),
            data_re_in(23) => data_re_in(1495),
            data_re_in(24) => data_re_in(1559),
            data_re_in(25) => data_re_in(1623),
            data_re_in(26) => data_re_in(1687),
            data_re_in(27) => data_re_in(1751),
            data_re_in(28) => data_re_in(1815),
            data_re_in(29) => data_re_in(1879),
            data_re_in(30) => data_re_in(1943),
            data_re_in(31) => data_re_in(2007),
            data_im_in(0) => data_im_in(23),
            data_im_in(1) => data_im_in(87),
            data_im_in(2) => data_im_in(151),
            data_im_in(3) => data_im_in(215),
            data_im_in(4) => data_im_in(279),
            data_im_in(5) => data_im_in(343),
            data_im_in(6) => data_im_in(407),
            data_im_in(7) => data_im_in(471),
            data_im_in(8) => data_im_in(535),
            data_im_in(9) => data_im_in(599),
            data_im_in(10) => data_im_in(663),
            data_im_in(11) => data_im_in(727),
            data_im_in(12) => data_im_in(791),
            data_im_in(13) => data_im_in(855),
            data_im_in(14) => data_im_in(919),
            data_im_in(15) => data_im_in(983),
            data_im_in(16) => data_im_in(1047),
            data_im_in(17) => data_im_in(1111),
            data_im_in(18) => data_im_in(1175),
            data_im_in(19) => data_im_in(1239),
            data_im_in(20) => data_im_in(1303),
            data_im_in(21) => data_im_in(1367),
            data_im_in(22) => data_im_in(1431),
            data_im_in(23) => data_im_in(1495),
            data_im_in(24) => data_im_in(1559),
            data_im_in(25) => data_im_in(1623),
            data_im_in(26) => data_im_in(1687),
            data_im_in(27) => data_im_in(1751),
            data_im_in(28) => data_im_in(1815),
            data_im_in(29) => data_im_in(1879),
            data_im_in(30) => data_im_in(1943),
            data_im_in(31) => data_im_in(2007),
            data_re_out(0) => first_stage_re_out(23),
            data_re_out(1) => first_stage_re_out(87),
            data_re_out(2) => first_stage_re_out(151),
            data_re_out(3) => first_stage_re_out(215),
            data_re_out(4) => first_stage_re_out(279),
            data_re_out(5) => first_stage_re_out(343),
            data_re_out(6) => first_stage_re_out(407),
            data_re_out(7) => first_stage_re_out(471),
            data_re_out(8) => first_stage_re_out(535),
            data_re_out(9) => first_stage_re_out(599),
            data_re_out(10) => first_stage_re_out(663),
            data_re_out(11) => first_stage_re_out(727),
            data_re_out(12) => first_stage_re_out(791),
            data_re_out(13) => first_stage_re_out(855),
            data_re_out(14) => first_stage_re_out(919),
            data_re_out(15) => first_stage_re_out(983),
            data_re_out(16) => first_stage_re_out(1047),
            data_re_out(17) => first_stage_re_out(1111),
            data_re_out(18) => first_stage_re_out(1175),
            data_re_out(19) => first_stage_re_out(1239),
            data_re_out(20) => first_stage_re_out(1303),
            data_re_out(21) => first_stage_re_out(1367),
            data_re_out(22) => first_stage_re_out(1431),
            data_re_out(23) => first_stage_re_out(1495),
            data_re_out(24) => first_stage_re_out(1559),
            data_re_out(25) => first_stage_re_out(1623),
            data_re_out(26) => first_stage_re_out(1687),
            data_re_out(27) => first_stage_re_out(1751),
            data_re_out(28) => first_stage_re_out(1815),
            data_re_out(29) => first_stage_re_out(1879),
            data_re_out(30) => first_stage_re_out(1943),
            data_re_out(31) => first_stage_re_out(2007),
            data_im_out(0) => first_stage_im_out(23),
            data_im_out(1) => first_stage_im_out(87),
            data_im_out(2) => first_stage_im_out(151),
            data_im_out(3) => first_stage_im_out(215),
            data_im_out(4) => first_stage_im_out(279),
            data_im_out(5) => first_stage_im_out(343),
            data_im_out(6) => first_stage_im_out(407),
            data_im_out(7) => first_stage_im_out(471),
            data_im_out(8) => first_stage_im_out(535),
            data_im_out(9) => first_stage_im_out(599),
            data_im_out(10) => first_stage_im_out(663),
            data_im_out(11) => first_stage_im_out(727),
            data_im_out(12) => first_stage_im_out(791),
            data_im_out(13) => first_stage_im_out(855),
            data_im_out(14) => first_stage_im_out(919),
            data_im_out(15) => first_stage_im_out(983),
            data_im_out(16) => first_stage_im_out(1047),
            data_im_out(17) => first_stage_im_out(1111),
            data_im_out(18) => first_stage_im_out(1175),
            data_im_out(19) => first_stage_im_out(1239),
            data_im_out(20) => first_stage_im_out(1303),
            data_im_out(21) => first_stage_im_out(1367),
            data_im_out(22) => first_stage_im_out(1431),
            data_im_out(23) => first_stage_im_out(1495),
            data_im_out(24) => first_stage_im_out(1559),
            data_im_out(25) => first_stage_im_out(1623),
            data_im_out(26) => first_stage_im_out(1687),
            data_im_out(27) => first_stage_im_out(1751),
            data_im_out(28) => first_stage_im_out(1815),
            data_im_out(29) => first_stage_im_out(1879),
            data_im_out(30) => first_stage_im_out(1943),
            data_im_out(31) => first_stage_im_out(2007)
        );

    ULFFT_PT32_24 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(24),
            data_re_in(1) => data_re_in(88),
            data_re_in(2) => data_re_in(152),
            data_re_in(3) => data_re_in(216),
            data_re_in(4) => data_re_in(280),
            data_re_in(5) => data_re_in(344),
            data_re_in(6) => data_re_in(408),
            data_re_in(7) => data_re_in(472),
            data_re_in(8) => data_re_in(536),
            data_re_in(9) => data_re_in(600),
            data_re_in(10) => data_re_in(664),
            data_re_in(11) => data_re_in(728),
            data_re_in(12) => data_re_in(792),
            data_re_in(13) => data_re_in(856),
            data_re_in(14) => data_re_in(920),
            data_re_in(15) => data_re_in(984),
            data_re_in(16) => data_re_in(1048),
            data_re_in(17) => data_re_in(1112),
            data_re_in(18) => data_re_in(1176),
            data_re_in(19) => data_re_in(1240),
            data_re_in(20) => data_re_in(1304),
            data_re_in(21) => data_re_in(1368),
            data_re_in(22) => data_re_in(1432),
            data_re_in(23) => data_re_in(1496),
            data_re_in(24) => data_re_in(1560),
            data_re_in(25) => data_re_in(1624),
            data_re_in(26) => data_re_in(1688),
            data_re_in(27) => data_re_in(1752),
            data_re_in(28) => data_re_in(1816),
            data_re_in(29) => data_re_in(1880),
            data_re_in(30) => data_re_in(1944),
            data_re_in(31) => data_re_in(2008),
            data_im_in(0) => data_im_in(24),
            data_im_in(1) => data_im_in(88),
            data_im_in(2) => data_im_in(152),
            data_im_in(3) => data_im_in(216),
            data_im_in(4) => data_im_in(280),
            data_im_in(5) => data_im_in(344),
            data_im_in(6) => data_im_in(408),
            data_im_in(7) => data_im_in(472),
            data_im_in(8) => data_im_in(536),
            data_im_in(9) => data_im_in(600),
            data_im_in(10) => data_im_in(664),
            data_im_in(11) => data_im_in(728),
            data_im_in(12) => data_im_in(792),
            data_im_in(13) => data_im_in(856),
            data_im_in(14) => data_im_in(920),
            data_im_in(15) => data_im_in(984),
            data_im_in(16) => data_im_in(1048),
            data_im_in(17) => data_im_in(1112),
            data_im_in(18) => data_im_in(1176),
            data_im_in(19) => data_im_in(1240),
            data_im_in(20) => data_im_in(1304),
            data_im_in(21) => data_im_in(1368),
            data_im_in(22) => data_im_in(1432),
            data_im_in(23) => data_im_in(1496),
            data_im_in(24) => data_im_in(1560),
            data_im_in(25) => data_im_in(1624),
            data_im_in(26) => data_im_in(1688),
            data_im_in(27) => data_im_in(1752),
            data_im_in(28) => data_im_in(1816),
            data_im_in(29) => data_im_in(1880),
            data_im_in(30) => data_im_in(1944),
            data_im_in(31) => data_im_in(2008),
            data_re_out(0) => first_stage_re_out(24),
            data_re_out(1) => first_stage_re_out(88),
            data_re_out(2) => first_stage_re_out(152),
            data_re_out(3) => first_stage_re_out(216),
            data_re_out(4) => first_stage_re_out(280),
            data_re_out(5) => first_stage_re_out(344),
            data_re_out(6) => first_stage_re_out(408),
            data_re_out(7) => first_stage_re_out(472),
            data_re_out(8) => first_stage_re_out(536),
            data_re_out(9) => first_stage_re_out(600),
            data_re_out(10) => first_stage_re_out(664),
            data_re_out(11) => first_stage_re_out(728),
            data_re_out(12) => first_stage_re_out(792),
            data_re_out(13) => first_stage_re_out(856),
            data_re_out(14) => first_stage_re_out(920),
            data_re_out(15) => first_stage_re_out(984),
            data_re_out(16) => first_stage_re_out(1048),
            data_re_out(17) => first_stage_re_out(1112),
            data_re_out(18) => first_stage_re_out(1176),
            data_re_out(19) => first_stage_re_out(1240),
            data_re_out(20) => first_stage_re_out(1304),
            data_re_out(21) => first_stage_re_out(1368),
            data_re_out(22) => first_stage_re_out(1432),
            data_re_out(23) => first_stage_re_out(1496),
            data_re_out(24) => first_stage_re_out(1560),
            data_re_out(25) => first_stage_re_out(1624),
            data_re_out(26) => first_stage_re_out(1688),
            data_re_out(27) => first_stage_re_out(1752),
            data_re_out(28) => first_stage_re_out(1816),
            data_re_out(29) => first_stage_re_out(1880),
            data_re_out(30) => first_stage_re_out(1944),
            data_re_out(31) => first_stage_re_out(2008),
            data_im_out(0) => first_stage_im_out(24),
            data_im_out(1) => first_stage_im_out(88),
            data_im_out(2) => first_stage_im_out(152),
            data_im_out(3) => first_stage_im_out(216),
            data_im_out(4) => first_stage_im_out(280),
            data_im_out(5) => first_stage_im_out(344),
            data_im_out(6) => first_stage_im_out(408),
            data_im_out(7) => first_stage_im_out(472),
            data_im_out(8) => first_stage_im_out(536),
            data_im_out(9) => first_stage_im_out(600),
            data_im_out(10) => first_stage_im_out(664),
            data_im_out(11) => first_stage_im_out(728),
            data_im_out(12) => first_stage_im_out(792),
            data_im_out(13) => first_stage_im_out(856),
            data_im_out(14) => first_stage_im_out(920),
            data_im_out(15) => first_stage_im_out(984),
            data_im_out(16) => first_stage_im_out(1048),
            data_im_out(17) => first_stage_im_out(1112),
            data_im_out(18) => first_stage_im_out(1176),
            data_im_out(19) => first_stage_im_out(1240),
            data_im_out(20) => first_stage_im_out(1304),
            data_im_out(21) => first_stage_im_out(1368),
            data_im_out(22) => first_stage_im_out(1432),
            data_im_out(23) => first_stage_im_out(1496),
            data_im_out(24) => first_stage_im_out(1560),
            data_im_out(25) => first_stage_im_out(1624),
            data_im_out(26) => first_stage_im_out(1688),
            data_im_out(27) => first_stage_im_out(1752),
            data_im_out(28) => first_stage_im_out(1816),
            data_im_out(29) => first_stage_im_out(1880),
            data_im_out(30) => first_stage_im_out(1944),
            data_im_out(31) => first_stage_im_out(2008)
        );

    ULFFT_PT32_25 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(25),
            data_re_in(1) => data_re_in(89),
            data_re_in(2) => data_re_in(153),
            data_re_in(3) => data_re_in(217),
            data_re_in(4) => data_re_in(281),
            data_re_in(5) => data_re_in(345),
            data_re_in(6) => data_re_in(409),
            data_re_in(7) => data_re_in(473),
            data_re_in(8) => data_re_in(537),
            data_re_in(9) => data_re_in(601),
            data_re_in(10) => data_re_in(665),
            data_re_in(11) => data_re_in(729),
            data_re_in(12) => data_re_in(793),
            data_re_in(13) => data_re_in(857),
            data_re_in(14) => data_re_in(921),
            data_re_in(15) => data_re_in(985),
            data_re_in(16) => data_re_in(1049),
            data_re_in(17) => data_re_in(1113),
            data_re_in(18) => data_re_in(1177),
            data_re_in(19) => data_re_in(1241),
            data_re_in(20) => data_re_in(1305),
            data_re_in(21) => data_re_in(1369),
            data_re_in(22) => data_re_in(1433),
            data_re_in(23) => data_re_in(1497),
            data_re_in(24) => data_re_in(1561),
            data_re_in(25) => data_re_in(1625),
            data_re_in(26) => data_re_in(1689),
            data_re_in(27) => data_re_in(1753),
            data_re_in(28) => data_re_in(1817),
            data_re_in(29) => data_re_in(1881),
            data_re_in(30) => data_re_in(1945),
            data_re_in(31) => data_re_in(2009),
            data_im_in(0) => data_im_in(25),
            data_im_in(1) => data_im_in(89),
            data_im_in(2) => data_im_in(153),
            data_im_in(3) => data_im_in(217),
            data_im_in(4) => data_im_in(281),
            data_im_in(5) => data_im_in(345),
            data_im_in(6) => data_im_in(409),
            data_im_in(7) => data_im_in(473),
            data_im_in(8) => data_im_in(537),
            data_im_in(9) => data_im_in(601),
            data_im_in(10) => data_im_in(665),
            data_im_in(11) => data_im_in(729),
            data_im_in(12) => data_im_in(793),
            data_im_in(13) => data_im_in(857),
            data_im_in(14) => data_im_in(921),
            data_im_in(15) => data_im_in(985),
            data_im_in(16) => data_im_in(1049),
            data_im_in(17) => data_im_in(1113),
            data_im_in(18) => data_im_in(1177),
            data_im_in(19) => data_im_in(1241),
            data_im_in(20) => data_im_in(1305),
            data_im_in(21) => data_im_in(1369),
            data_im_in(22) => data_im_in(1433),
            data_im_in(23) => data_im_in(1497),
            data_im_in(24) => data_im_in(1561),
            data_im_in(25) => data_im_in(1625),
            data_im_in(26) => data_im_in(1689),
            data_im_in(27) => data_im_in(1753),
            data_im_in(28) => data_im_in(1817),
            data_im_in(29) => data_im_in(1881),
            data_im_in(30) => data_im_in(1945),
            data_im_in(31) => data_im_in(2009),
            data_re_out(0) => first_stage_re_out(25),
            data_re_out(1) => first_stage_re_out(89),
            data_re_out(2) => first_stage_re_out(153),
            data_re_out(3) => first_stage_re_out(217),
            data_re_out(4) => first_stage_re_out(281),
            data_re_out(5) => first_stage_re_out(345),
            data_re_out(6) => first_stage_re_out(409),
            data_re_out(7) => first_stage_re_out(473),
            data_re_out(8) => first_stage_re_out(537),
            data_re_out(9) => first_stage_re_out(601),
            data_re_out(10) => first_stage_re_out(665),
            data_re_out(11) => first_stage_re_out(729),
            data_re_out(12) => first_stage_re_out(793),
            data_re_out(13) => first_stage_re_out(857),
            data_re_out(14) => first_stage_re_out(921),
            data_re_out(15) => first_stage_re_out(985),
            data_re_out(16) => first_stage_re_out(1049),
            data_re_out(17) => first_stage_re_out(1113),
            data_re_out(18) => first_stage_re_out(1177),
            data_re_out(19) => first_stage_re_out(1241),
            data_re_out(20) => first_stage_re_out(1305),
            data_re_out(21) => first_stage_re_out(1369),
            data_re_out(22) => first_stage_re_out(1433),
            data_re_out(23) => first_stage_re_out(1497),
            data_re_out(24) => first_stage_re_out(1561),
            data_re_out(25) => first_stage_re_out(1625),
            data_re_out(26) => first_stage_re_out(1689),
            data_re_out(27) => first_stage_re_out(1753),
            data_re_out(28) => first_stage_re_out(1817),
            data_re_out(29) => first_stage_re_out(1881),
            data_re_out(30) => first_stage_re_out(1945),
            data_re_out(31) => first_stage_re_out(2009),
            data_im_out(0) => first_stage_im_out(25),
            data_im_out(1) => first_stage_im_out(89),
            data_im_out(2) => first_stage_im_out(153),
            data_im_out(3) => first_stage_im_out(217),
            data_im_out(4) => first_stage_im_out(281),
            data_im_out(5) => first_stage_im_out(345),
            data_im_out(6) => first_stage_im_out(409),
            data_im_out(7) => first_stage_im_out(473),
            data_im_out(8) => first_stage_im_out(537),
            data_im_out(9) => first_stage_im_out(601),
            data_im_out(10) => first_stage_im_out(665),
            data_im_out(11) => first_stage_im_out(729),
            data_im_out(12) => first_stage_im_out(793),
            data_im_out(13) => first_stage_im_out(857),
            data_im_out(14) => first_stage_im_out(921),
            data_im_out(15) => first_stage_im_out(985),
            data_im_out(16) => first_stage_im_out(1049),
            data_im_out(17) => first_stage_im_out(1113),
            data_im_out(18) => first_stage_im_out(1177),
            data_im_out(19) => first_stage_im_out(1241),
            data_im_out(20) => first_stage_im_out(1305),
            data_im_out(21) => first_stage_im_out(1369),
            data_im_out(22) => first_stage_im_out(1433),
            data_im_out(23) => first_stage_im_out(1497),
            data_im_out(24) => first_stage_im_out(1561),
            data_im_out(25) => first_stage_im_out(1625),
            data_im_out(26) => first_stage_im_out(1689),
            data_im_out(27) => first_stage_im_out(1753),
            data_im_out(28) => first_stage_im_out(1817),
            data_im_out(29) => first_stage_im_out(1881),
            data_im_out(30) => first_stage_im_out(1945),
            data_im_out(31) => first_stage_im_out(2009)
        );

    ULFFT_PT32_26 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(26),
            data_re_in(1) => data_re_in(90),
            data_re_in(2) => data_re_in(154),
            data_re_in(3) => data_re_in(218),
            data_re_in(4) => data_re_in(282),
            data_re_in(5) => data_re_in(346),
            data_re_in(6) => data_re_in(410),
            data_re_in(7) => data_re_in(474),
            data_re_in(8) => data_re_in(538),
            data_re_in(9) => data_re_in(602),
            data_re_in(10) => data_re_in(666),
            data_re_in(11) => data_re_in(730),
            data_re_in(12) => data_re_in(794),
            data_re_in(13) => data_re_in(858),
            data_re_in(14) => data_re_in(922),
            data_re_in(15) => data_re_in(986),
            data_re_in(16) => data_re_in(1050),
            data_re_in(17) => data_re_in(1114),
            data_re_in(18) => data_re_in(1178),
            data_re_in(19) => data_re_in(1242),
            data_re_in(20) => data_re_in(1306),
            data_re_in(21) => data_re_in(1370),
            data_re_in(22) => data_re_in(1434),
            data_re_in(23) => data_re_in(1498),
            data_re_in(24) => data_re_in(1562),
            data_re_in(25) => data_re_in(1626),
            data_re_in(26) => data_re_in(1690),
            data_re_in(27) => data_re_in(1754),
            data_re_in(28) => data_re_in(1818),
            data_re_in(29) => data_re_in(1882),
            data_re_in(30) => data_re_in(1946),
            data_re_in(31) => data_re_in(2010),
            data_im_in(0) => data_im_in(26),
            data_im_in(1) => data_im_in(90),
            data_im_in(2) => data_im_in(154),
            data_im_in(3) => data_im_in(218),
            data_im_in(4) => data_im_in(282),
            data_im_in(5) => data_im_in(346),
            data_im_in(6) => data_im_in(410),
            data_im_in(7) => data_im_in(474),
            data_im_in(8) => data_im_in(538),
            data_im_in(9) => data_im_in(602),
            data_im_in(10) => data_im_in(666),
            data_im_in(11) => data_im_in(730),
            data_im_in(12) => data_im_in(794),
            data_im_in(13) => data_im_in(858),
            data_im_in(14) => data_im_in(922),
            data_im_in(15) => data_im_in(986),
            data_im_in(16) => data_im_in(1050),
            data_im_in(17) => data_im_in(1114),
            data_im_in(18) => data_im_in(1178),
            data_im_in(19) => data_im_in(1242),
            data_im_in(20) => data_im_in(1306),
            data_im_in(21) => data_im_in(1370),
            data_im_in(22) => data_im_in(1434),
            data_im_in(23) => data_im_in(1498),
            data_im_in(24) => data_im_in(1562),
            data_im_in(25) => data_im_in(1626),
            data_im_in(26) => data_im_in(1690),
            data_im_in(27) => data_im_in(1754),
            data_im_in(28) => data_im_in(1818),
            data_im_in(29) => data_im_in(1882),
            data_im_in(30) => data_im_in(1946),
            data_im_in(31) => data_im_in(2010),
            data_re_out(0) => first_stage_re_out(26),
            data_re_out(1) => first_stage_re_out(90),
            data_re_out(2) => first_stage_re_out(154),
            data_re_out(3) => first_stage_re_out(218),
            data_re_out(4) => first_stage_re_out(282),
            data_re_out(5) => first_stage_re_out(346),
            data_re_out(6) => first_stage_re_out(410),
            data_re_out(7) => first_stage_re_out(474),
            data_re_out(8) => first_stage_re_out(538),
            data_re_out(9) => first_stage_re_out(602),
            data_re_out(10) => first_stage_re_out(666),
            data_re_out(11) => first_stage_re_out(730),
            data_re_out(12) => first_stage_re_out(794),
            data_re_out(13) => first_stage_re_out(858),
            data_re_out(14) => first_stage_re_out(922),
            data_re_out(15) => first_stage_re_out(986),
            data_re_out(16) => first_stage_re_out(1050),
            data_re_out(17) => first_stage_re_out(1114),
            data_re_out(18) => first_stage_re_out(1178),
            data_re_out(19) => first_stage_re_out(1242),
            data_re_out(20) => first_stage_re_out(1306),
            data_re_out(21) => first_stage_re_out(1370),
            data_re_out(22) => first_stage_re_out(1434),
            data_re_out(23) => first_stage_re_out(1498),
            data_re_out(24) => first_stage_re_out(1562),
            data_re_out(25) => first_stage_re_out(1626),
            data_re_out(26) => first_stage_re_out(1690),
            data_re_out(27) => first_stage_re_out(1754),
            data_re_out(28) => first_stage_re_out(1818),
            data_re_out(29) => first_stage_re_out(1882),
            data_re_out(30) => first_stage_re_out(1946),
            data_re_out(31) => first_stage_re_out(2010),
            data_im_out(0) => first_stage_im_out(26),
            data_im_out(1) => first_stage_im_out(90),
            data_im_out(2) => first_stage_im_out(154),
            data_im_out(3) => first_stage_im_out(218),
            data_im_out(4) => first_stage_im_out(282),
            data_im_out(5) => first_stage_im_out(346),
            data_im_out(6) => first_stage_im_out(410),
            data_im_out(7) => first_stage_im_out(474),
            data_im_out(8) => first_stage_im_out(538),
            data_im_out(9) => first_stage_im_out(602),
            data_im_out(10) => first_stage_im_out(666),
            data_im_out(11) => first_stage_im_out(730),
            data_im_out(12) => first_stage_im_out(794),
            data_im_out(13) => first_stage_im_out(858),
            data_im_out(14) => first_stage_im_out(922),
            data_im_out(15) => first_stage_im_out(986),
            data_im_out(16) => first_stage_im_out(1050),
            data_im_out(17) => first_stage_im_out(1114),
            data_im_out(18) => first_stage_im_out(1178),
            data_im_out(19) => first_stage_im_out(1242),
            data_im_out(20) => first_stage_im_out(1306),
            data_im_out(21) => first_stage_im_out(1370),
            data_im_out(22) => first_stage_im_out(1434),
            data_im_out(23) => first_stage_im_out(1498),
            data_im_out(24) => first_stage_im_out(1562),
            data_im_out(25) => first_stage_im_out(1626),
            data_im_out(26) => first_stage_im_out(1690),
            data_im_out(27) => first_stage_im_out(1754),
            data_im_out(28) => first_stage_im_out(1818),
            data_im_out(29) => first_stage_im_out(1882),
            data_im_out(30) => first_stage_im_out(1946),
            data_im_out(31) => first_stage_im_out(2010)
        );

    ULFFT_PT32_27 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(27),
            data_re_in(1) => data_re_in(91),
            data_re_in(2) => data_re_in(155),
            data_re_in(3) => data_re_in(219),
            data_re_in(4) => data_re_in(283),
            data_re_in(5) => data_re_in(347),
            data_re_in(6) => data_re_in(411),
            data_re_in(7) => data_re_in(475),
            data_re_in(8) => data_re_in(539),
            data_re_in(9) => data_re_in(603),
            data_re_in(10) => data_re_in(667),
            data_re_in(11) => data_re_in(731),
            data_re_in(12) => data_re_in(795),
            data_re_in(13) => data_re_in(859),
            data_re_in(14) => data_re_in(923),
            data_re_in(15) => data_re_in(987),
            data_re_in(16) => data_re_in(1051),
            data_re_in(17) => data_re_in(1115),
            data_re_in(18) => data_re_in(1179),
            data_re_in(19) => data_re_in(1243),
            data_re_in(20) => data_re_in(1307),
            data_re_in(21) => data_re_in(1371),
            data_re_in(22) => data_re_in(1435),
            data_re_in(23) => data_re_in(1499),
            data_re_in(24) => data_re_in(1563),
            data_re_in(25) => data_re_in(1627),
            data_re_in(26) => data_re_in(1691),
            data_re_in(27) => data_re_in(1755),
            data_re_in(28) => data_re_in(1819),
            data_re_in(29) => data_re_in(1883),
            data_re_in(30) => data_re_in(1947),
            data_re_in(31) => data_re_in(2011),
            data_im_in(0) => data_im_in(27),
            data_im_in(1) => data_im_in(91),
            data_im_in(2) => data_im_in(155),
            data_im_in(3) => data_im_in(219),
            data_im_in(4) => data_im_in(283),
            data_im_in(5) => data_im_in(347),
            data_im_in(6) => data_im_in(411),
            data_im_in(7) => data_im_in(475),
            data_im_in(8) => data_im_in(539),
            data_im_in(9) => data_im_in(603),
            data_im_in(10) => data_im_in(667),
            data_im_in(11) => data_im_in(731),
            data_im_in(12) => data_im_in(795),
            data_im_in(13) => data_im_in(859),
            data_im_in(14) => data_im_in(923),
            data_im_in(15) => data_im_in(987),
            data_im_in(16) => data_im_in(1051),
            data_im_in(17) => data_im_in(1115),
            data_im_in(18) => data_im_in(1179),
            data_im_in(19) => data_im_in(1243),
            data_im_in(20) => data_im_in(1307),
            data_im_in(21) => data_im_in(1371),
            data_im_in(22) => data_im_in(1435),
            data_im_in(23) => data_im_in(1499),
            data_im_in(24) => data_im_in(1563),
            data_im_in(25) => data_im_in(1627),
            data_im_in(26) => data_im_in(1691),
            data_im_in(27) => data_im_in(1755),
            data_im_in(28) => data_im_in(1819),
            data_im_in(29) => data_im_in(1883),
            data_im_in(30) => data_im_in(1947),
            data_im_in(31) => data_im_in(2011),
            data_re_out(0) => first_stage_re_out(27),
            data_re_out(1) => first_stage_re_out(91),
            data_re_out(2) => first_stage_re_out(155),
            data_re_out(3) => first_stage_re_out(219),
            data_re_out(4) => first_stage_re_out(283),
            data_re_out(5) => first_stage_re_out(347),
            data_re_out(6) => first_stage_re_out(411),
            data_re_out(7) => first_stage_re_out(475),
            data_re_out(8) => first_stage_re_out(539),
            data_re_out(9) => first_stage_re_out(603),
            data_re_out(10) => first_stage_re_out(667),
            data_re_out(11) => first_stage_re_out(731),
            data_re_out(12) => first_stage_re_out(795),
            data_re_out(13) => first_stage_re_out(859),
            data_re_out(14) => first_stage_re_out(923),
            data_re_out(15) => first_stage_re_out(987),
            data_re_out(16) => first_stage_re_out(1051),
            data_re_out(17) => first_stage_re_out(1115),
            data_re_out(18) => first_stage_re_out(1179),
            data_re_out(19) => first_stage_re_out(1243),
            data_re_out(20) => first_stage_re_out(1307),
            data_re_out(21) => first_stage_re_out(1371),
            data_re_out(22) => first_stage_re_out(1435),
            data_re_out(23) => first_stage_re_out(1499),
            data_re_out(24) => first_stage_re_out(1563),
            data_re_out(25) => first_stage_re_out(1627),
            data_re_out(26) => first_stage_re_out(1691),
            data_re_out(27) => first_stage_re_out(1755),
            data_re_out(28) => first_stage_re_out(1819),
            data_re_out(29) => first_stage_re_out(1883),
            data_re_out(30) => first_stage_re_out(1947),
            data_re_out(31) => first_stage_re_out(2011),
            data_im_out(0) => first_stage_im_out(27),
            data_im_out(1) => first_stage_im_out(91),
            data_im_out(2) => first_stage_im_out(155),
            data_im_out(3) => first_stage_im_out(219),
            data_im_out(4) => first_stage_im_out(283),
            data_im_out(5) => first_stage_im_out(347),
            data_im_out(6) => first_stage_im_out(411),
            data_im_out(7) => first_stage_im_out(475),
            data_im_out(8) => first_stage_im_out(539),
            data_im_out(9) => first_stage_im_out(603),
            data_im_out(10) => first_stage_im_out(667),
            data_im_out(11) => first_stage_im_out(731),
            data_im_out(12) => first_stage_im_out(795),
            data_im_out(13) => first_stage_im_out(859),
            data_im_out(14) => first_stage_im_out(923),
            data_im_out(15) => first_stage_im_out(987),
            data_im_out(16) => first_stage_im_out(1051),
            data_im_out(17) => first_stage_im_out(1115),
            data_im_out(18) => first_stage_im_out(1179),
            data_im_out(19) => first_stage_im_out(1243),
            data_im_out(20) => first_stage_im_out(1307),
            data_im_out(21) => first_stage_im_out(1371),
            data_im_out(22) => first_stage_im_out(1435),
            data_im_out(23) => first_stage_im_out(1499),
            data_im_out(24) => first_stage_im_out(1563),
            data_im_out(25) => first_stage_im_out(1627),
            data_im_out(26) => first_stage_im_out(1691),
            data_im_out(27) => first_stage_im_out(1755),
            data_im_out(28) => first_stage_im_out(1819),
            data_im_out(29) => first_stage_im_out(1883),
            data_im_out(30) => first_stage_im_out(1947),
            data_im_out(31) => first_stage_im_out(2011)
        );

    ULFFT_PT32_28 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(28),
            data_re_in(1) => data_re_in(92),
            data_re_in(2) => data_re_in(156),
            data_re_in(3) => data_re_in(220),
            data_re_in(4) => data_re_in(284),
            data_re_in(5) => data_re_in(348),
            data_re_in(6) => data_re_in(412),
            data_re_in(7) => data_re_in(476),
            data_re_in(8) => data_re_in(540),
            data_re_in(9) => data_re_in(604),
            data_re_in(10) => data_re_in(668),
            data_re_in(11) => data_re_in(732),
            data_re_in(12) => data_re_in(796),
            data_re_in(13) => data_re_in(860),
            data_re_in(14) => data_re_in(924),
            data_re_in(15) => data_re_in(988),
            data_re_in(16) => data_re_in(1052),
            data_re_in(17) => data_re_in(1116),
            data_re_in(18) => data_re_in(1180),
            data_re_in(19) => data_re_in(1244),
            data_re_in(20) => data_re_in(1308),
            data_re_in(21) => data_re_in(1372),
            data_re_in(22) => data_re_in(1436),
            data_re_in(23) => data_re_in(1500),
            data_re_in(24) => data_re_in(1564),
            data_re_in(25) => data_re_in(1628),
            data_re_in(26) => data_re_in(1692),
            data_re_in(27) => data_re_in(1756),
            data_re_in(28) => data_re_in(1820),
            data_re_in(29) => data_re_in(1884),
            data_re_in(30) => data_re_in(1948),
            data_re_in(31) => data_re_in(2012),
            data_im_in(0) => data_im_in(28),
            data_im_in(1) => data_im_in(92),
            data_im_in(2) => data_im_in(156),
            data_im_in(3) => data_im_in(220),
            data_im_in(4) => data_im_in(284),
            data_im_in(5) => data_im_in(348),
            data_im_in(6) => data_im_in(412),
            data_im_in(7) => data_im_in(476),
            data_im_in(8) => data_im_in(540),
            data_im_in(9) => data_im_in(604),
            data_im_in(10) => data_im_in(668),
            data_im_in(11) => data_im_in(732),
            data_im_in(12) => data_im_in(796),
            data_im_in(13) => data_im_in(860),
            data_im_in(14) => data_im_in(924),
            data_im_in(15) => data_im_in(988),
            data_im_in(16) => data_im_in(1052),
            data_im_in(17) => data_im_in(1116),
            data_im_in(18) => data_im_in(1180),
            data_im_in(19) => data_im_in(1244),
            data_im_in(20) => data_im_in(1308),
            data_im_in(21) => data_im_in(1372),
            data_im_in(22) => data_im_in(1436),
            data_im_in(23) => data_im_in(1500),
            data_im_in(24) => data_im_in(1564),
            data_im_in(25) => data_im_in(1628),
            data_im_in(26) => data_im_in(1692),
            data_im_in(27) => data_im_in(1756),
            data_im_in(28) => data_im_in(1820),
            data_im_in(29) => data_im_in(1884),
            data_im_in(30) => data_im_in(1948),
            data_im_in(31) => data_im_in(2012),
            data_re_out(0) => first_stage_re_out(28),
            data_re_out(1) => first_stage_re_out(92),
            data_re_out(2) => first_stage_re_out(156),
            data_re_out(3) => first_stage_re_out(220),
            data_re_out(4) => first_stage_re_out(284),
            data_re_out(5) => first_stage_re_out(348),
            data_re_out(6) => first_stage_re_out(412),
            data_re_out(7) => first_stage_re_out(476),
            data_re_out(8) => first_stage_re_out(540),
            data_re_out(9) => first_stage_re_out(604),
            data_re_out(10) => first_stage_re_out(668),
            data_re_out(11) => first_stage_re_out(732),
            data_re_out(12) => first_stage_re_out(796),
            data_re_out(13) => first_stage_re_out(860),
            data_re_out(14) => first_stage_re_out(924),
            data_re_out(15) => first_stage_re_out(988),
            data_re_out(16) => first_stage_re_out(1052),
            data_re_out(17) => first_stage_re_out(1116),
            data_re_out(18) => first_stage_re_out(1180),
            data_re_out(19) => first_stage_re_out(1244),
            data_re_out(20) => first_stage_re_out(1308),
            data_re_out(21) => first_stage_re_out(1372),
            data_re_out(22) => first_stage_re_out(1436),
            data_re_out(23) => first_stage_re_out(1500),
            data_re_out(24) => first_stage_re_out(1564),
            data_re_out(25) => first_stage_re_out(1628),
            data_re_out(26) => first_stage_re_out(1692),
            data_re_out(27) => first_stage_re_out(1756),
            data_re_out(28) => first_stage_re_out(1820),
            data_re_out(29) => first_stage_re_out(1884),
            data_re_out(30) => first_stage_re_out(1948),
            data_re_out(31) => first_stage_re_out(2012),
            data_im_out(0) => first_stage_im_out(28),
            data_im_out(1) => first_stage_im_out(92),
            data_im_out(2) => first_stage_im_out(156),
            data_im_out(3) => first_stage_im_out(220),
            data_im_out(4) => first_stage_im_out(284),
            data_im_out(5) => first_stage_im_out(348),
            data_im_out(6) => first_stage_im_out(412),
            data_im_out(7) => first_stage_im_out(476),
            data_im_out(8) => first_stage_im_out(540),
            data_im_out(9) => first_stage_im_out(604),
            data_im_out(10) => first_stage_im_out(668),
            data_im_out(11) => first_stage_im_out(732),
            data_im_out(12) => first_stage_im_out(796),
            data_im_out(13) => first_stage_im_out(860),
            data_im_out(14) => first_stage_im_out(924),
            data_im_out(15) => first_stage_im_out(988),
            data_im_out(16) => first_stage_im_out(1052),
            data_im_out(17) => first_stage_im_out(1116),
            data_im_out(18) => first_stage_im_out(1180),
            data_im_out(19) => first_stage_im_out(1244),
            data_im_out(20) => first_stage_im_out(1308),
            data_im_out(21) => first_stage_im_out(1372),
            data_im_out(22) => first_stage_im_out(1436),
            data_im_out(23) => first_stage_im_out(1500),
            data_im_out(24) => first_stage_im_out(1564),
            data_im_out(25) => first_stage_im_out(1628),
            data_im_out(26) => first_stage_im_out(1692),
            data_im_out(27) => first_stage_im_out(1756),
            data_im_out(28) => first_stage_im_out(1820),
            data_im_out(29) => first_stage_im_out(1884),
            data_im_out(30) => first_stage_im_out(1948),
            data_im_out(31) => first_stage_im_out(2012)
        );

    ULFFT_PT32_29 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(29),
            data_re_in(1) => data_re_in(93),
            data_re_in(2) => data_re_in(157),
            data_re_in(3) => data_re_in(221),
            data_re_in(4) => data_re_in(285),
            data_re_in(5) => data_re_in(349),
            data_re_in(6) => data_re_in(413),
            data_re_in(7) => data_re_in(477),
            data_re_in(8) => data_re_in(541),
            data_re_in(9) => data_re_in(605),
            data_re_in(10) => data_re_in(669),
            data_re_in(11) => data_re_in(733),
            data_re_in(12) => data_re_in(797),
            data_re_in(13) => data_re_in(861),
            data_re_in(14) => data_re_in(925),
            data_re_in(15) => data_re_in(989),
            data_re_in(16) => data_re_in(1053),
            data_re_in(17) => data_re_in(1117),
            data_re_in(18) => data_re_in(1181),
            data_re_in(19) => data_re_in(1245),
            data_re_in(20) => data_re_in(1309),
            data_re_in(21) => data_re_in(1373),
            data_re_in(22) => data_re_in(1437),
            data_re_in(23) => data_re_in(1501),
            data_re_in(24) => data_re_in(1565),
            data_re_in(25) => data_re_in(1629),
            data_re_in(26) => data_re_in(1693),
            data_re_in(27) => data_re_in(1757),
            data_re_in(28) => data_re_in(1821),
            data_re_in(29) => data_re_in(1885),
            data_re_in(30) => data_re_in(1949),
            data_re_in(31) => data_re_in(2013),
            data_im_in(0) => data_im_in(29),
            data_im_in(1) => data_im_in(93),
            data_im_in(2) => data_im_in(157),
            data_im_in(3) => data_im_in(221),
            data_im_in(4) => data_im_in(285),
            data_im_in(5) => data_im_in(349),
            data_im_in(6) => data_im_in(413),
            data_im_in(7) => data_im_in(477),
            data_im_in(8) => data_im_in(541),
            data_im_in(9) => data_im_in(605),
            data_im_in(10) => data_im_in(669),
            data_im_in(11) => data_im_in(733),
            data_im_in(12) => data_im_in(797),
            data_im_in(13) => data_im_in(861),
            data_im_in(14) => data_im_in(925),
            data_im_in(15) => data_im_in(989),
            data_im_in(16) => data_im_in(1053),
            data_im_in(17) => data_im_in(1117),
            data_im_in(18) => data_im_in(1181),
            data_im_in(19) => data_im_in(1245),
            data_im_in(20) => data_im_in(1309),
            data_im_in(21) => data_im_in(1373),
            data_im_in(22) => data_im_in(1437),
            data_im_in(23) => data_im_in(1501),
            data_im_in(24) => data_im_in(1565),
            data_im_in(25) => data_im_in(1629),
            data_im_in(26) => data_im_in(1693),
            data_im_in(27) => data_im_in(1757),
            data_im_in(28) => data_im_in(1821),
            data_im_in(29) => data_im_in(1885),
            data_im_in(30) => data_im_in(1949),
            data_im_in(31) => data_im_in(2013),
            data_re_out(0) => first_stage_re_out(29),
            data_re_out(1) => first_stage_re_out(93),
            data_re_out(2) => first_stage_re_out(157),
            data_re_out(3) => first_stage_re_out(221),
            data_re_out(4) => first_stage_re_out(285),
            data_re_out(5) => first_stage_re_out(349),
            data_re_out(6) => first_stage_re_out(413),
            data_re_out(7) => first_stage_re_out(477),
            data_re_out(8) => first_stage_re_out(541),
            data_re_out(9) => first_stage_re_out(605),
            data_re_out(10) => first_stage_re_out(669),
            data_re_out(11) => first_stage_re_out(733),
            data_re_out(12) => first_stage_re_out(797),
            data_re_out(13) => first_stage_re_out(861),
            data_re_out(14) => first_stage_re_out(925),
            data_re_out(15) => first_stage_re_out(989),
            data_re_out(16) => first_stage_re_out(1053),
            data_re_out(17) => first_stage_re_out(1117),
            data_re_out(18) => first_stage_re_out(1181),
            data_re_out(19) => first_stage_re_out(1245),
            data_re_out(20) => first_stage_re_out(1309),
            data_re_out(21) => first_stage_re_out(1373),
            data_re_out(22) => first_stage_re_out(1437),
            data_re_out(23) => first_stage_re_out(1501),
            data_re_out(24) => first_stage_re_out(1565),
            data_re_out(25) => first_stage_re_out(1629),
            data_re_out(26) => first_stage_re_out(1693),
            data_re_out(27) => first_stage_re_out(1757),
            data_re_out(28) => first_stage_re_out(1821),
            data_re_out(29) => first_stage_re_out(1885),
            data_re_out(30) => first_stage_re_out(1949),
            data_re_out(31) => first_stage_re_out(2013),
            data_im_out(0) => first_stage_im_out(29),
            data_im_out(1) => first_stage_im_out(93),
            data_im_out(2) => first_stage_im_out(157),
            data_im_out(3) => first_stage_im_out(221),
            data_im_out(4) => first_stage_im_out(285),
            data_im_out(5) => first_stage_im_out(349),
            data_im_out(6) => first_stage_im_out(413),
            data_im_out(7) => first_stage_im_out(477),
            data_im_out(8) => first_stage_im_out(541),
            data_im_out(9) => first_stage_im_out(605),
            data_im_out(10) => first_stage_im_out(669),
            data_im_out(11) => first_stage_im_out(733),
            data_im_out(12) => first_stage_im_out(797),
            data_im_out(13) => first_stage_im_out(861),
            data_im_out(14) => first_stage_im_out(925),
            data_im_out(15) => first_stage_im_out(989),
            data_im_out(16) => first_stage_im_out(1053),
            data_im_out(17) => first_stage_im_out(1117),
            data_im_out(18) => first_stage_im_out(1181),
            data_im_out(19) => first_stage_im_out(1245),
            data_im_out(20) => first_stage_im_out(1309),
            data_im_out(21) => first_stage_im_out(1373),
            data_im_out(22) => first_stage_im_out(1437),
            data_im_out(23) => first_stage_im_out(1501),
            data_im_out(24) => first_stage_im_out(1565),
            data_im_out(25) => first_stage_im_out(1629),
            data_im_out(26) => first_stage_im_out(1693),
            data_im_out(27) => first_stage_im_out(1757),
            data_im_out(28) => first_stage_im_out(1821),
            data_im_out(29) => first_stage_im_out(1885),
            data_im_out(30) => first_stage_im_out(1949),
            data_im_out(31) => first_stage_im_out(2013)
        );

    ULFFT_PT32_30 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(30),
            data_re_in(1) => data_re_in(94),
            data_re_in(2) => data_re_in(158),
            data_re_in(3) => data_re_in(222),
            data_re_in(4) => data_re_in(286),
            data_re_in(5) => data_re_in(350),
            data_re_in(6) => data_re_in(414),
            data_re_in(7) => data_re_in(478),
            data_re_in(8) => data_re_in(542),
            data_re_in(9) => data_re_in(606),
            data_re_in(10) => data_re_in(670),
            data_re_in(11) => data_re_in(734),
            data_re_in(12) => data_re_in(798),
            data_re_in(13) => data_re_in(862),
            data_re_in(14) => data_re_in(926),
            data_re_in(15) => data_re_in(990),
            data_re_in(16) => data_re_in(1054),
            data_re_in(17) => data_re_in(1118),
            data_re_in(18) => data_re_in(1182),
            data_re_in(19) => data_re_in(1246),
            data_re_in(20) => data_re_in(1310),
            data_re_in(21) => data_re_in(1374),
            data_re_in(22) => data_re_in(1438),
            data_re_in(23) => data_re_in(1502),
            data_re_in(24) => data_re_in(1566),
            data_re_in(25) => data_re_in(1630),
            data_re_in(26) => data_re_in(1694),
            data_re_in(27) => data_re_in(1758),
            data_re_in(28) => data_re_in(1822),
            data_re_in(29) => data_re_in(1886),
            data_re_in(30) => data_re_in(1950),
            data_re_in(31) => data_re_in(2014),
            data_im_in(0) => data_im_in(30),
            data_im_in(1) => data_im_in(94),
            data_im_in(2) => data_im_in(158),
            data_im_in(3) => data_im_in(222),
            data_im_in(4) => data_im_in(286),
            data_im_in(5) => data_im_in(350),
            data_im_in(6) => data_im_in(414),
            data_im_in(7) => data_im_in(478),
            data_im_in(8) => data_im_in(542),
            data_im_in(9) => data_im_in(606),
            data_im_in(10) => data_im_in(670),
            data_im_in(11) => data_im_in(734),
            data_im_in(12) => data_im_in(798),
            data_im_in(13) => data_im_in(862),
            data_im_in(14) => data_im_in(926),
            data_im_in(15) => data_im_in(990),
            data_im_in(16) => data_im_in(1054),
            data_im_in(17) => data_im_in(1118),
            data_im_in(18) => data_im_in(1182),
            data_im_in(19) => data_im_in(1246),
            data_im_in(20) => data_im_in(1310),
            data_im_in(21) => data_im_in(1374),
            data_im_in(22) => data_im_in(1438),
            data_im_in(23) => data_im_in(1502),
            data_im_in(24) => data_im_in(1566),
            data_im_in(25) => data_im_in(1630),
            data_im_in(26) => data_im_in(1694),
            data_im_in(27) => data_im_in(1758),
            data_im_in(28) => data_im_in(1822),
            data_im_in(29) => data_im_in(1886),
            data_im_in(30) => data_im_in(1950),
            data_im_in(31) => data_im_in(2014),
            data_re_out(0) => first_stage_re_out(30),
            data_re_out(1) => first_stage_re_out(94),
            data_re_out(2) => first_stage_re_out(158),
            data_re_out(3) => first_stage_re_out(222),
            data_re_out(4) => first_stage_re_out(286),
            data_re_out(5) => first_stage_re_out(350),
            data_re_out(6) => first_stage_re_out(414),
            data_re_out(7) => first_stage_re_out(478),
            data_re_out(8) => first_stage_re_out(542),
            data_re_out(9) => first_stage_re_out(606),
            data_re_out(10) => first_stage_re_out(670),
            data_re_out(11) => first_stage_re_out(734),
            data_re_out(12) => first_stage_re_out(798),
            data_re_out(13) => first_stage_re_out(862),
            data_re_out(14) => first_stage_re_out(926),
            data_re_out(15) => first_stage_re_out(990),
            data_re_out(16) => first_stage_re_out(1054),
            data_re_out(17) => first_stage_re_out(1118),
            data_re_out(18) => first_stage_re_out(1182),
            data_re_out(19) => first_stage_re_out(1246),
            data_re_out(20) => first_stage_re_out(1310),
            data_re_out(21) => first_stage_re_out(1374),
            data_re_out(22) => first_stage_re_out(1438),
            data_re_out(23) => first_stage_re_out(1502),
            data_re_out(24) => first_stage_re_out(1566),
            data_re_out(25) => first_stage_re_out(1630),
            data_re_out(26) => first_stage_re_out(1694),
            data_re_out(27) => first_stage_re_out(1758),
            data_re_out(28) => first_stage_re_out(1822),
            data_re_out(29) => first_stage_re_out(1886),
            data_re_out(30) => first_stage_re_out(1950),
            data_re_out(31) => first_stage_re_out(2014),
            data_im_out(0) => first_stage_im_out(30),
            data_im_out(1) => first_stage_im_out(94),
            data_im_out(2) => first_stage_im_out(158),
            data_im_out(3) => first_stage_im_out(222),
            data_im_out(4) => first_stage_im_out(286),
            data_im_out(5) => first_stage_im_out(350),
            data_im_out(6) => first_stage_im_out(414),
            data_im_out(7) => first_stage_im_out(478),
            data_im_out(8) => first_stage_im_out(542),
            data_im_out(9) => first_stage_im_out(606),
            data_im_out(10) => first_stage_im_out(670),
            data_im_out(11) => first_stage_im_out(734),
            data_im_out(12) => first_stage_im_out(798),
            data_im_out(13) => first_stage_im_out(862),
            data_im_out(14) => first_stage_im_out(926),
            data_im_out(15) => first_stage_im_out(990),
            data_im_out(16) => first_stage_im_out(1054),
            data_im_out(17) => first_stage_im_out(1118),
            data_im_out(18) => first_stage_im_out(1182),
            data_im_out(19) => first_stage_im_out(1246),
            data_im_out(20) => first_stage_im_out(1310),
            data_im_out(21) => first_stage_im_out(1374),
            data_im_out(22) => first_stage_im_out(1438),
            data_im_out(23) => first_stage_im_out(1502),
            data_im_out(24) => first_stage_im_out(1566),
            data_im_out(25) => first_stage_im_out(1630),
            data_im_out(26) => first_stage_im_out(1694),
            data_im_out(27) => first_stage_im_out(1758),
            data_im_out(28) => first_stage_im_out(1822),
            data_im_out(29) => first_stage_im_out(1886),
            data_im_out(30) => first_stage_im_out(1950),
            data_im_out(31) => first_stage_im_out(2014)
        );

    ULFFT_PT32_31 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(31),
            data_re_in(1) => data_re_in(95),
            data_re_in(2) => data_re_in(159),
            data_re_in(3) => data_re_in(223),
            data_re_in(4) => data_re_in(287),
            data_re_in(5) => data_re_in(351),
            data_re_in(6) => data_re_in(415),
            data_re_in(7) => data_re_in(479),
            data_re_in(8) => data_re_in(543),
            data_re_in(9) => data_re_in(607),
            data_re_in(10) => data_re_in(671),
            data_re_in(11) => data_re_in(735),
            data_re_in(12) => data_re_in(799),
            data_re_in(13) => data_re_in(863),
            data_re_in(14) => data_re_in(927),
            data_re_in(15) => data_re_in(991),
            data_re_in(16) => data_re_in(1055),
            data_re_in(17) => data_re_in(1119),
            data_re_in(18) => data_re_in(1183),
            data_re_in(19) => data_re_in(1247),
            data_re_in(20) => data_re_in(1311),
            data_re_in(21) => data_re_in(1375),
            data_re_in(22) => data_re_in(1439),
            data_re_in(23) => data_re_in(1503),
            data_re_in(24) => data_re_in(1567),
            data_re_in(25) => data_re_in(1631),
            data_re_in(26) => data_re_in(1695),
            data_re_in(27) => data_re_in(1759),
            data_re_in(28) => data_re_in(1823),
            data_re_in(29) => data_re_in(1887),
            data_re_in(30) => data_re_in(1951),
            data_re_in(31) => data_re_in(2015),
            data_im_in(0) => data_im_in(31),
            data_im_in(1) => data_im_in(95),
            data_im_in(2) => data_im_in(159),
            data_im_in(3) => data_im_in(223),
            data_im_in(4) => data_im_in(287),
            data_im_in(5) => data_im_in(351),
            data_im_in(6) => data_im_in(415),
            data_im_in(7) => data_im_in(479),
            data_im_in(8) => data_im_in(543),
            data_im_in(9) => data_im_in(607),
            data_im_in(10) => data_im_in(671),
            data_im_in(11) => data_im_in(735),
            data_im_in(12) => data_im_in(799),
            data_im_in(13) => data_im_in(863),
            data_im_in(14) => data_im_in(927),
            data_im_in(15) => data_im_in(991),
            data_im_in(16) => data_im_in(1055),
            data_im_in(17) => data_im_in(1119),
            data_im_in(18) => data_im_in(1183),
            data_im_in(19) => data_im_in(1247),
            data_im_in(20) => data_im_in(1311),
            data_im_in(21) => data_im_in(1375),
            data_im_in(22) => data_im_in(1439),
            data_im_in(23) => data_im_in(1503),
            data_im_in(24) => data_im_in(1567),
            data_im_in(25) => data_im_in(1631),
            data_im_in(26) => data_im_in(1695),
            data_im_in(27) => data_im_in(1759),
            data_im_in(28) => data_im_in(1823),
            data_im_in(29) => data_im_in(1887),
            data_im_in(30) => data_im_in(1951),
            data_im_in(31) => data_im_in(2015),
            data_re_out(0) => first_stage_re_out(31),
            data_re_out(1) => first_stage_re_out(95),
            data_re_out(2) => first_stage_re_out(159),
            data_re_out(3) => first_stage_re_out(223),
            data_re_out(4) => first_stage_re_out(287),
            data_re_out(5) => first_stage_re_out(351),
            data_re_out(6) => first_stage_re_out(415),
            data_re_out(7) => first_stage_re_out(479),
            data_re_out(8) => first_stage_re_out(543),
            data_re_out(9) => first_stage_re_out(607),
            data_re_out(10) => first_stage_re_out(671),
            data_re_out(11) => first_stage_re_out(735),
            data_re_out(12) => first_stage_re_out(799),
            data_re_out(13) => first_stage_re_out(863),
            data_re_out(14) => first_stage_re_out(927),
            data_re_out(15) => first_stage_re_out(991),
            data_re_out(16) => first_stage_re_out(1055),
            data_re_out(17) => first_stage_re_out(1119),
            data_re_out(18) => first_stage_re_out(1183),
            data_re_out(19) => first_stage_re_out(1247),
            data_re_out(20) => first_stage_re_out(1311),
            data_re_out(21) => first_stage_re_out(1375),
            data_re_out(22) => first_stage_re_out(1439),
            data_re_out(23) => first_stage_re_out(1503),
            data_re_out(24) => first_stage_re_out(1567),
            data_re_out(25) => first_stage_re_out(1631),
            data_re_out(26) => first_stage_re_out(1695),
            data_re_out(27) => first_stage_re_out(1759),
            data_re_out(28) => first_stage_re_out(1823),
            data_re_out(29) => first_stage_re_out(1887),
            data_re_out(30) => first_stage_re_out(1951),
            data_re_out(31) => first_stage_re_out(2015),
            data_im_out(0) => first_stage_im_out(31),
            data_im_out(1) => first_stage_im_out(95),
            data_im_out(2) => first_stage_im_out(159),
            data_im_out(3) => first_stage_im_out(223),
            data_im_out(4) => first_stage_im_out(287),
            data_im_out(5) => first_stage_im_out(351),
            data_im_out(6) => first_stage_im_out(415),
            data_im_out(7) => first_stage_im_out(479),
            data_im_out(8) => first_stage_im_out(543),
            data_im_out(9) => first_stage_im_out(607),
            data_im_out(10) => first_stage_im_out(671),
            data_im_out(11) => first_stage_im_out(735),
            data_im_out(12) => first_stage_im_out(799),
            data_im_out(13) => first_stage_im_out(863),
            data_im_out(14) => first_stage_im_out(927),
            data_im_out(15) => first_stage_im_out(991),
            data_im_out(16) => first_stage_im_out(1055),
            data_im_out(17) => first_stage_im_out(1119),
            data_im_out(18) => first_stage_im_out(1183),
            data_im_out(19) => first_stage_im_out(1247),
            data_im_out(20) => first_stage_im_out(1311),
            data_im_out(21) => first_stage_im_out(1375),
            data_im_out(22) => first_stage_im_out(1439),
            data_im_out(23) => first_stage_im_out(1503),
            data_im_out(24) => first_stage_im_out(1567),
            data_im_out(25) => first_stage_im_out(1631),
            data_im_out(26) => first_stage_im_out(1695),
            data_im_out(27) => first_stage_im_out(1759),
            data_im_out(28) => first_stage_im_out(1823),
            data_im_out(29) => first_stage_im_out(1887),
            data_im_out(30) => first_stage_im_out(1951),
            data_im_out(31) => first_stage_im_out(2015)
        );

    ULFFT_PT32_32 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(32),
            data_re_in(1) => data_re_in(96),
            data_re_in(2) => data_re_in(160),
            data_re_in(3) => data_re_in(224),
            data_re_in(4) => data_re_in(288),
            data_re_in(5) => data_re_in(352),
            data_re_in(6) => data_re_in(416),
            data_re_in(7) => data_re_in(480),
            data_re_in(8) => data_re_in(544),
            data_re_in(9) => data_re_in(608),
            data_re_in(10) => data_re_in(672),
            data_re_in(11) => data_re_in(736),
            data_re_in(12) => data_re_in(800),
            data_re_in(13) => data_re_in(864),
            data_re_in(14) => data_re_in(928),
            data_re_in(15) => data_re_in(992),
            data_re_in(16) => data_re_in(1056),
            data_re_in(17) => data_re_in(1120),
            data_re_in(18) => data_re_in(1184),
            data_re_in(19) => data_re_in(1248),
            data_re_in(20) => data_re_in(1312),
            data_re_in(21) => data_re_in(1376),
            data_re_in(22) => data_re_in(1440),
            data_re_in(23) => data_re_in(1504),
            data_re_in(24) => data_re_in(1568),
            data_re_in(25) => data_re_in(1632),
            data_re_in(26) => data_re_in(1696),
            data_re_in(27) => data_re_in(1760),
            data_re_in(28) => data_re_in(1824),
            data_re_in(29) => data_re_in(1888),
            data_re_in(30) => data_re_in(1952),
            data_re_in(31) => data_re_in(2016),
            data_im_in(0) => data_im_in(32),
            data_im_in(1) => data_im_in(96),
            data_im_in(2) => data_im_in(160),
            data_im_in(3) => data_im_in(224),
            data_im_in(4) => data_im_in(288),
            data_im_in(5) => data_im_in(352),
            data_im_in(6) => data_im_in(416),
            data_im_in(7) => data_im_in(480),
            data_im_in(8) => data_im_in(544),
            data_im_in(9) => data_im_in(608),
            data_im_in(10) => data_im_in(672),
            data_im_in(11) => data_im_in(736),
            data_im_in(12) => data_im_in(800),
            data_im_in(13) => data_im_in(864),
            data_im_in(14) => data_im_in(928),
            data_im_in(15) => data_im_in(992),
            data_im_in(16) => data_im_in(1056),
            data_im_in(17) => data_im_in(1120),
            data_im_in(18) => data_im_in(1184),
            data_im_in(19) => data_im_in(1248),
            data_im_in(20) => data_im_in(1312),
            data_im_in(21) => data_im_in(1376),
            data_im_in(22) => data_im_in(1440),
            data_im_in(23) => data_im_in(1504),
            data_im_in(24) => data_im_in(1568),
            data_im_in(25) => data_im_in(1632),
            data_im_in(26) => data_im_in(1696),
            data_im_in(27) => data_im_in(1760),
            data_im_in(28) => data_im_in(1824),
            data_im_in(29) => data_im_in(1888),
            data_im_in(30) => data_im_in(1952),
            data_im_in(31) => data_im_in(2016),
            data_re_out(0) => first_stage_re_out(32),
            data_re_out(1) => first_stage_re_out(96),
            data_re_out(2) => first_stage_re_out(160),
            data_re_out(3) => first_stage_re_out(224),
            data_re_out(4) => first_stage_re_out(288),
            data_re_out(5) => first_stage_re_out(352),
            data_re_out(6) => first_stage_re_out(416),
            data_re_out(7) => first_stage_re_out(480),
            data_re_out(8) => first_stage_re_out(544),
            data_re_out(9) => first_stage_re_out(608),
            data_re_out(10) => first_stage_re_out(672),
            data_re_out(11) => first_stage_re_out(736),
            data_re_out(12) => first_stage_re_out(800),
            data_re_out(13) => first_stage_re_out(864),
            data_re_out(14) => first_stage_re_out(928),
            data_re_out(15) => first_stage_re_out(992),
            data_re_out(16) => first_stage_re_out(1056),
            data_re_out(17) => first_stage_re_out(1120),
            data_re_out(18) => first_stage_re_out(1184),
            data_re_out(19) => first_stage_re_out(1248),
            data_re_out(20) => first_stage_re_out(1312),
            data_re_out(21) => first_stage_re_out(1376),
            data_re_out(22) => first_stage_re_out(1440),
            data_re_out(23) => first_stage_re_out(1504),
            data_re_out(24) => first_stage_re_out(1568),
            data_re_out(25) => first_stage_re_out(1632),
            data_re_out(26) => first_stage_re_out(1696),
            data_re_out(27) => first_stage_re_out(1760),
            data_re_out(28) => first_stage_re_out(1824),
            data_re_out(29) => first_stage_re_out(1888),
            data_re_out(30) => first_stage_re_out(1952),
            data_re_out(31) => first_stage_re_out(2016),
            data_im_out(0) => first_stage_im_out(32),
            data_im_out(1) => first_stage_im_out(96),
            data_im_out(2) => first_stage_im_out(160),
            data_im_out(3) => first_stage_im_out(224),
            data_im_out(4) => first_stage_im_out(288),
            data_im_out(5) => first_stage_im_out(352),
            data_im_out(6) => first_stage_im_out(416),
            data_im_out(7) => first_stage_im_out(480),
            data_im_out(8) => first_stage_im_out(544),
            data_im_out(9) => first_stage_im_out(608),
            data_im_out(10) => first_stage_im_out(672),
            data_im_out(11) => first_stage_im_out(736),
            data_im_out(12) => first_stage_im_out(800),
            data_im_out(13) => first_stage_im_out(864),
            data_im_out(14) => first_stage_im_out(928),
            data_im_out(15) => first_stage_im_out(992),
            data_im_out(16) => first_stage_im_out(1056),
            data_im_out(17) => first_stage_im_out(1120),
            data_im_out(18) => first_stage_im_out(1184),
            data_im_out(19) => first_stage_im_out(1248),
            data_im_out(20) => first_stage_im_out(1312),
            data_im_out(21) => first_stage_im_out(1376),
            data_im_out(22) => first_stage_im_out(1440),
            data_im_out(23) => first_stage_im_out(1504),
            data_im_out(24) => first_stage_im_out(1568),
            data_im_out(25) => first_stage_im_out(1632),
            data_im_out(26) => first_stage_im_out(1696),
            data_im_out(27) => first_stage_im_out(1760),
            data_im_out(28) => first_stage_im_out(1824),
            data_im_out(29) => first_stage_im_out(1888),
            data_im_out(30) => first_stage_im_out(1952),
            data_im_out(31) => first_stage_im_out(2016)
        );

    ULFFT_PT32_33 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(33),
            data_re_in(1) => data_re_in(97),
            data_re_in(2) => data_re_in(161),
            data_re_in(3) => data_re_in(225),
            data_re_in(4) => data_re_in(289),
            data_re_in(5) => data_re_in(353),
            data_re_in(6) => data_re_in(417),
            data_re_in(7) => data_re_in(481),
            data_re_in(8) => data_re_in(545),
            data_re_in(9) => data_re_in(609),
            data_re_in(10) => data_re_in(673),
            data_re_in(11) => data_re_in(737),
            data_re_in(12) => data_re_in(801),
            data_re_in(13) => data_re_in(865),
            data_re_in(14) => data_re_in(929),
            data_re_in(15) => data_re_in(993),
            data_re_in(16) => data_re_in(1057),
            data_re_in(17) => data_re_in(1121),
            data_re_in(18) => data_re_in(1185),
            data_re_in(19) => data_re_in(1249),
            data_re_in(20) => data_re_in(1313),
            data_re_in(21) => data_re_in(1377),
            data_re_in(22) => data_re_in(1441),
            data_re_in(23) => data_re_in(1505),
            data_re_in(24) => data_re_in(1569),
            data_re_in(25) => data_re_in(1633),
            data_re_in(26) => data_re_in(1697),
            data_re_in(27) => data_re_in(1761),
            data_re_in(28) => data_re_in(1825),
            data_re_in(29) => data_re_in(1889),
            data_re_in(30) => data_re_in(1953),
            data_re_in(31) => data_re_in(2017),
            data_im_in(0) => data_im_in(33),
            data_im_in(1) => data_im_in(97),
            data_im_in(2) => data_im_in(161),
            data_im_in(3) => data_im_in(225),
            data_im_in(4) => data_im_in(289),
            data_im_in(5) => data_im_in(353),
            data_im_in(6) => data_im_in(417),
            data_im_in(7) => data_im_in(481),
            data_im_in(8) => data_im_in(545),
            data_im_in(9) => data_im_in(609),
            data_im_in(10) => data_im_in(673),
            data_im_in(11) => data_im_in(737),
            data_im_in(12) => data_im_in(801),
            data_im_in(13) => data_im_in(865),
            data_im_in(14) => data_im_in(929),
            data_im_in(15) => data_im_in(993),
            data_im_in(16) => data_im_in(1057),
            data_im_in(17) => data_im_in(1121),
            data_im_in(18) => data_im_in(1185),
            data_im_in(19) => data_im_in(1249),
            data_im_in(20) => data_im_in(1313),
            data_im_in(21) => data_im_in(1377),
            data_im_in(22) => data_im_in(1441),
            data_im_in(23) => data_im_in(1505),
            data_im_in(24) => data_im_in(1569),
            data_im_in(25) => data_im_in(1633),
            data_im_in(26) => data_im_in(1697),
            data_im_in(27) => data_im_in(1761),
            data_im_in(28) => data_im_in(1825),
            data_im_in(29) => data_im_in(1889),
            data_im_in(30) => data_im_in(1953),
            data_im_in(31) => data_im_in(2017),
            data_re_out(0) => first_stage_re_out(33),
            data_re_out(1) => first_stage_re_out(97),
            data_re_out(2) => first_stage_re_out(161),
            data_re_out(3) => first_stage_re_out(225),
            data_re_out(4) => first_stage_re_out(289),
            data_re_out(5) => first_stage_re_out(353),
            data_re_out(6) => first_stage_re_out(417),
            data_re_out(7) => first_stage_re_out(481),
            data_re_out(8) => first_stage_re_out(545),
            data_re_out(9) => first_stage_re_out(609),
            data_re_out(10) => first_stage_re_out(673),
            data_re_out(11) => first_stage_re_out(737),
            data_re_out(12) => first_stage_re_out(801),
            data_re_out(13) => first_stage_re_out(865),
            data_re_out(14) => first_stage_re_out(929),
            data_re_out(15) => first_stage_re_out(993),
            data_re_out(16) => first_stage_re_out(1057),
            data_re_out(17) => first_stage_re_out(1121),
            data_re_out(18) => first_stage_re_out(1185),
            data_re_out(19) => first_stage_re_out(1249),
            data_re_out(20) => first_stage_re_out(1313),
            data_re_out(21) => first_stage_re_out(1377),
            data_re_out(22) => first_stage_re_out(1441),
            data_re_out(23) => first_stage_re_out(1505),
            data_re_out(24) => first_stage_re_out(1569),
            data_re_out(25) => first_stage_re_out(1633),
            data_re_out(26) => first_stage_re_out(1697),
            data_re_out(27) => first_stage_re_out(1761),
            data_re_out(28) => first_stage_re_out(1825),
            data_re_out(29) => first_stage_re_out(1889),
            data_re_out(30) => first_stage_re_out(1953),
            data_re_out(31) => first_stage_re_out(2017),
            data_im_out(0) => first_stage_im_out(33),
            data_im_out(1) => first_stage_im_out(97),
            data_im_out(2) => first_stage_im_out(161),
            data_im_out(3) => first_stage_im_out(225),
            data_im_out(4) => first_stage_im_out(289),
            data_im_out(5) => first_stage_im_out(353),
            data_im_out(6) => first_stage_im_out(417),
            data_im_out(7) => first_stage_im_out(481),
            data_im_out(8) => first_stage_im_out(545),
            data_im_out(9) => first_stage_im_out(609),
            data_im_out(10) => first_stage_im_out(673),
            data_im_out(11) => first_stage_im_out(737),
            data_im_out(12) => first_stage_im_out(801),
            data_im_out(13) => first_stage_im_out(865),
            data_im_out(14) => first_stage_im_out(929),
            data_im_out(15) => first_stage_im_out(993),
            data_im_out(16) => first_stage_im_out(1057),
            data_im_out(17) => first_stage_im_out(1121),
            data_im_out(18) => first_stage_im_out(1185),
            data_im_out(19) => first_stage_im_out(1249),
            data_im_out(20) => first_stage_im_out(1313),
            data_im_out(21) => first_stage_im_out(1377),
            data_im_out(22) => first_stage_im_out(1441),
            data_im_out(23) => first_stage_im_out(1505),
            data_im_out(24) => first_stage_im_out(1569),
            data_im_out(25) => first_stage_im_out(1633),
            data_im_out(26) => first_stage_im_out(1697),
            data_im_out(27) => first_stage_im_out(1761),
            data_im_out(28) => first_stage_im_out(1825),
            data_im_out(29) => first_stage_im_out(1889),
            data_im_out(30) => first_stage_im_out(1953),
            data_im_out(31) => first_stage_im_out(2017)
        );

    ULFFT_PT32_34 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(34),
            data_re_in(1) => data_re_in(98),
            data_re_in(2) => data_re_in(162),
            data_re_in(3) => data_re_in(226),
            data_re_in(4) => data_re_in(290),
            data_re_in(5) => data_re_in(354),
            data_re_in(6) => data_re_in(418),
            data_re_in(7) => data_re_in(482),
            data_re_in(8) => data_re_in(546),
            data_re_in(9) => data_re_in(610),
            data_re_in(10) => data_re_in(674),
            data_re_in(11) => data_re_in(738),
            data_re_in(12) => data_re_in(802),
            data_re_in(13) => data_re_in(866),
            data_re_in(14) => data_re_in(930),
            data_re_in(15) => data_re_in(994),
            data_re_in(16) => data_re_in(1058),
            data_re_in(17) => data_re_in(1122),
            data_re_in(18) => data_re_in(1186),
            data_re_in(19) => data_re_in(1250),
            data_re_in(20) => data_re_in(1314),
            data_re_in(21) => data_re_in(1378),
            data_re_in(22) => data_re_in(1442),
            data_re_in(23) => data_re_in(1506),
            data_re_in(24) => data_re_in(1570),
            data_re_in(25) => data_re_in(1634),
            data_re_in(26) => data_re_in(1698),
            data_re_in(27) => data_re_in(1762),
            data_re_in(28) => data_re_in(1826),
            data_re_in(29) => data_re_in(1890),
            data_re_in(30) => data_re_in(1954),
            data_re_in(31) => data_re_in(2018),
            data_im_in(0) => data_im_in(34),
            data_im_in(1) => data_im_in(98),
            data_im_in(2) => data_im_in(162),
            data_im_in(3) => data_im_in(226),
            data_im_in(4) => data_im_in(290),
            data_im_in(5) => data_im_in(354),
            data_im_in(6) => data_im_in(418),
            data_im_in(7) => data_im_in(482),
            data_im_in(8) => data_im_in(546),
            data_im_in(9) => data_im_in(610),
            data_im_in(10) => data_im_in(674),
            data_im_in(11) => data_im_in(738),
            data_im_in(12) => data_im_in(802),
            data_im_in(13) => data_im_in(866),
            data_im_in(14) => data_im_in(930),
            data_im_in(15) => data_im_in(994),
            data_im_in(16) => data_im_in(1058),
            data_im_in(17) => data_im_in(1122),
            data_im_in(18) => data_im_in(1186),
            data_im_in(19) => data_im_in(1250),
            data_im_in(20) => data_im_in(1314),
            data_im_in(21) => data_im_in(1378),
            data_im_in(22) => data_im_in(1442),
            data_im_in(23) => data_im_in(1506),
            data_im_in(24) => data_im_in(1570),
            data_im_in(25) => data_im_in(1634),
            data_im_in(26) => data_im_in(1698),
            data_im_in(27) => data_im_in(1762),
            data_im_in(28) => data_im_in(1826),
            data_im_in(29) => data_im_in(1890),
            data_im_in(30) => data_im_in(1954),
            data_im_in(31) => data_im_in(2018),
            data_re_out(0) => first_stage_re_out(34),
            data_re_out(1) => first_stage_re_out(98),
            data_re_out(2) => first_stage_re_out(162),
            data_re_out(3) => first_stage_re_out(226),
            data_re_out(4) => first_stage_re_out(290),
            data_re_out(5) => first_stage_re_out(354),
            data_re_out(6) => first_stage_re_out(418),
            data_re_out(7) => first_stage_re_out(482),
            data_re_out(8) => first_stage_re_out(546),
            data_re_out(9) => first_stage_re_out(610),
            data_re_out(10) => first_stage_re_out(674),
            data_re_out(11) => first_stage_re_out(738),
            data_re_out(12) => first_stage_re_out(802),
            data_re_out(13) => first_stage_re_out(866),
            data_re_out(14) => first_stage_re_out(930),
            data_re_out(15) => first_stage_re_out(994),
            data_re_out(16) => first_stage_re_out(1058),
            data_re_out(17) => first_stage_re_out(1122),
            data_re_out(18) => first_stage_re_out(1186),
            data_re_out(19) => first_stage_re_out(1250),
            data_re_out(20) => first_stage_re_out(1314),
            data_re_out(21) => first_stage_re_out(1378),
            data_re_out(22) => first_stage_re_out(1442),
            data_re_out(23) => first_stage_re_out(1506),
            data_re_out(24) => first_stage_re_out(1570),
            data_re_out(25) => first_stage_re_out(1634),
            data_re_out(26) => first_stage_re_out(1698),
            data_re_out(27) => first_stage_re_out(1762),
            data_re_out(28) => first_stage_re_out(1826),
            data_re_out(29) => first_stage_re_out(1890),
            data_re_out(30) => first_stage_re_out(1954),
            data_re_out(31) => first_stage_re_out(2018),
            data_im_out(0) => first_stage_im_out(34),
            data_im_out(1) => first_stage_im_out(98),
            data_im_out(2) => first_stage_im_out(162),
            data_im_out(3) => first_stage_im_out(226),
            data_im_out(4) => first_stage_im_out(290),
            data_im_out(5) => first_stage_im_out(354),
            data_im_out(6) => first_stage_im_out(418),
            data_im_out(7) => first_stage_im_out(482),
            data_im_out(8) => first_stage_im_out(546),
            data_im_out(9) => first_stage_im_out(610),
            data_im_out(10) => first_stage_im_out(674),
            data_im_out(11) => first_stage_im_out(738),
            data_im_out(12) => first_stage_im_out(802),
            data_im_out(13) => first_stage_im_out(866),
            data_im_out(14) => first_stage_im_out(930),
            data_im_out(15) => first_stage_im_out(994),
            data_im_out(16) => first_stage_im_out(1058),
            data_im_out(17) => first_stage_im_out(1122),
            data_im_out(18) => first_stage_im_out(1186),
            data_im_out(19) => first_stage_im_out(1250),
            data_im_out(20) => first_stage_im_out(1314),
            data_im_out(21) => first_stage_im_out(1378),
            data_im_out(22) => first_stage_im_out(1442),
            data_im_out(23) => first_stage_im_out(1506),
            data_im_out(24) => first_stage_im_out(1570),
            data_im_out(25) => first_stage_im_out(1634),
            data_im_out(26) => first_stage_im_out(1698),
            data_im_out(27) => first_stage_im_out(1762),
            data_im_out(28) => first_stage_im_out(1826),
            data_im_out(29) => first_stage_im_out(1890),
            data_im_out(30) => first_stage_im_out(1954),
            data_im_out(31) => first_stage_im_out(2018)
        );

    ULFFT_PT32_35 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(35),
            data_re_in(1) => data_re_in(99),
            data_re_in(2) => data_re_in(163),
            data_re_in(3) => data_re_in(227),
            data_re_in(4) => data_re_in(291),
            data_re_in(5) => data_re_in(355),
            data_re_in(6) => data_re_in(419),
            data_re_in(7) => data_re_in(483),
            data_re_in(8) => data_re_in(547),
            data_re_in(9) => data_re_in(611),
            data_re_in(10) => data_re_in(675),
            data_re_in(11) => data_re_in(739),
            data_re_in(12) => data_re_in(803),
            data_re_in(13) => data_re_in(867),
            data_re_in(14) => data_re_in(931),
            data_re_in(15) => data_re_in(995),
            data_re_in(16) => data_re_in(1059),
            data_re_in(17) => data_re_in(1123),
            data_re_in(18) => data_re_in(1187),
            data_re_in(19) => data_re_in(1251),
            data_re_in(20) => data_re_in(1315),
            data_re_in(21) => data_re_in(1379),
            data_re_in(22) => data_re_in(1443),
            data_re_in(23) => data_re_in(1507),
            data_re_in(24) => data_re_in(1571),
            data_re_in(25) => data_re_in(1635),
            data_re_in(26) => data_re_in(1699),
            data_re_in(27) => data_re_in(1763),
            data_re_in(28) => data_re_in(1827),
            data_re_in(29) => data_re_in(1891),
            data_re_in(30) => data_re_in(1955),
            data_re_in(31) => data_re_in(2019),
            data_im_in(0) => data_im_in(35),
            data_im_in(1) => data_im_in(99),
            data_im_in(2) => data_im_in(163),
            data_im_in(3) => data_im_in(227),
            data_im_in(4) => data_im_in(291),
            data_im_in(5) => data_im_in(355),
            data_im_in(6) => data_im_in(419),
            data_im_in(7) => data_im_in(483),
            data_im_in(8) => data_im_in(547),
            data_im_in(9) => data_im_in(611),
            data_im_in(10) => data_im_in(675),
            data_im_in(11) => data_im_in(739),
            data_im_in(12) => data_im_in(803),
            data_im_in(13) => data_im_in(867),
            data_im_in(14) => data_im_in(931),
            data_im_in(15) => data_im_in(995),
            data_im_in(16) => data_im_in(1059),
            data_im_in(17) => data_im_in(1123),
            data_im_in(18) => data_im_in(1187),
            data_im_in(19) => data_im_in(1251),
            data_im_in(20) => data_im_in(1315),
            data_im_in(21) => data_im_in(1379),
            data_im_in(22) => data_im_in(1443),
            data_im_in(23) => data_im_in(1507),
            data_im_in(24) => data_im_in(1571),
            data_im_in(25) => data_im_in(1635),
            data_im_in(26) => data_im_in(1699),
            data_im_in(27) => data_im_in(1763),
            data_im_in(28) => data_im_in(1827),
            data_im_in(29) => data_im_in(1891),
            data_im_in(30) => data_im_in(1955),
            data_im_in(31) => data_im_in(2019),
            data_re_out(0) => first_stage_re_out(35),
            data_re_out(1) => first_stage_re_out(99),
            data_re_out(2) => first_stage_re_out(163),
            data_re_out(3) => first_stage_re_out(227),
            data_re_out(4) => first_stage_re_out(291),
            data_re_out(5) => first_stage_re_out(355),
            data_re_out(6) => first_stage_re_out(419),
            data_re_out(7) => first_stage_re_out(483),
            data_re_out(8) => first_stage_re_out(547),
            data_re_out(9) => first_stage_re_out(611),
            data_re_out(10) => first_stage_re_out(675),
            data_re_out(11) => first_stage_re_out(739),
            data_re_out(12) => first_stage_re_out(803),
            data_re_out(13) => first_stage_re_out(867),
            data_re_out(14) => first_stage_re_out(931),
            data_re_out(15) => first_stage_re_out(995),
            data_re_out(16) => first_stage_re_out(1059),
            data_re_out(17) => first_stage_re_out(1123),
            data_re_out(18) => first_stage_re_out(1187),
            data_re_out(19) => first_stage_re_out(1251),
            data_re_out(20) => first_stage_re_out(1315),
            data_re_out(21) => first_stage_re_out(1379),
            data_re_out(22) => first_stage_re_out(1443),
            data_re_out(23) => first_stage_re_out(1507),
            data_re_out(24) => first_stage_re_out(1571),
            data_re_out(25) => first_stage_re_out(1635),
            data_re_out(26) => first_stage_re_out(1699),
            data_re_out(27) => first_stage_re_out(1763),
            data_re_out(28) => first_stage_re_out(1827),
            data_re_out(29) => first_stage_re_out(1891),
            data_re_out(30) => first_stage_re_out(1955),
            data_re_out(31) => first_stage_re_out(2019),
            data_im_out(0) => first_stage_im_out(35),
            data_im_out(1) => first_stage_im_out(99),
            data_im_out(2) => first_stage_im_out(163),
            data_im_out(3) => first_stage_im_out(227),
            data_im_out(4) => first_stage_im_out(291),
            data_im_out(5) => first_stage_im_out(355),
            data_im_out(6) => first_stage_im_out(419),
            data_im_out(7) => first_stage_im_out(483),
            data_im_out(8) => first_stage_im_out(547),
            data_im_out(9) => first_stage_im_out(611),
            data_im_out(10) => first_stage_im_out(675),
            data_im_out(11) => first_stage_im_out(739),
            data_im_out(12) => first_stage_im_out(803),
            data_im_out(13) => first_stage_im_out(867),
            data_im_out(14) => first_stage_im_out(931),
            data_im_out(15) => first_stage_im_out(995),
            data_im_out(16) => first_stage_im_out(1059),
            data_im_out(17) => first_stage_im_out(1123),
            data_im_out(18) => first_stage_im_out(1187),
            data_im_out(19) => first_stage_im_out(1251),
            data_im_out(20) => first_stage_im_out(1315),
            data_im_out(21) => first_stage_im_out(1379),
            data_im_out(22) => first_stage_im_out(1443),
            data_im_out(23) => first_stage_im_out(1507),
            data_im_out(24) => first_stage_im_out(1571),
            data_im_out(25) => first_stage_im_out(1635),
            data_im_out(26) => first_stage_im_out(1699),
            data_im_out(27) => first_stage_im_out(1763),
            data_im_out(28) => first_stage_im_out(1827),
            data_im_out(29) => first_stage_im_out(1891),
            data_im_out(30) => first_stage_im_out(1955),
            data_im_out(31) => first_stage_im_out(2019)
        );

    ULFFT_PT32_36 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(36),
            data_re_in(1) => data_re_in(100),
            data_re_in(2) => data_re_in(164),
            data_re_in(3) => data_re_in(228),
            data_re_in(4) => data_re_in(292),
            data_re_in(5) => data_re_in(356),
            data_re_in(6) => data_re_in(420),
            data_re_in(7) => data_re_in(484),
            data_re_in(8) => data_re_in(548),
            data_re_in(9) => data_re_in(612),
            data_re_in(10) => data_re_in(676),
            data_re_in(11) => data_re_in(740),
            data_re_in(12) => data_re_in(804),
            data_re_in(13) => data_re_in(868),
            data_re_in(14) => data_re_in(932),
            data_re_in(15) => data_re_in(996),
            data_re_in(16) => data_re_in(1060),
            data_re_in(17) => data_re_in(1124),
            data_re_in(18) => data_re_in(1188),
            data_re_in(19) => data_re_in(1252),
            data_re_in(20) => data_re_in(1316),
            data_re_in(21) => data_re_in(1380),
            data_re_in(22) => data_re_in(1444),
            data_re_in(23) => data_re_in(1508),
            data_re_in(24) => data_re_in(1572),
            data_re_in(25) => data_re_in(1636),
            data_re_in(26) => data_re_in(1700),
            data_re_in(27) => data_re_in(1764),
            data_re_in(28) => data_re_in(1828),
            data_re_in(29) => data_re_in(1892),
            data_re_in(30) => data_re_in(1956),
            data_re_in(31) => data_re_in(2020),
            data_im_in(0) => data_im_in(36),
            data_im_in(1) => data_im_in(100),
            data_im_in(2) => data_im_in(164),
            data_im_in(3) => data_im_in(228),
            data_im_in(4) => data_im_in(292),
            data_im_in(5) => data_im_in(356),
            data_im_in(6) => data_im_in(420),
            data_im_in(7) => data_im_in(484),
            data_im_in(8) => data_im_in(548),
            data_im_in(9) => data_im_in(612),
            data_im_in(10) => data_im_in(676),
            data_im_in(11) => data_im_in(740),
            data_im_in(12) => data_im_in(804),
            data_im_in(13) => data_im_in(868),
            data_im_in(14) => data_im_in(932),
            data_im_in(15) => data_im_in(996),
            data_im_in(16) => data_im_in(1060),
            data_im_in(17) => data_im_in(1124),
            data_im_in(18) => data_im_in(1188),
            data_im_in(19) => data_im_in(1252),
            data_im_in(20) => data_im_in(1316),
            data_im_in(21) => data_im_in(1380),
            data_im_in(22) => data_im_in(1444),
            data_im_in(23) => data_im_in(1508),
            data_im_in(24) => data_im_in(1572),
            data_im_in(25) => data_im_in(1636),
            data_im_in(26) => data_im_in(1700),
            data_im_in(27) => data_im_in(1764),
            data_im_in(28) => data_im_in(1828),
            data_im_in(29) => data_im_in(1892),
            data_im_in(30) => data_im_in(1956),
            data_im_in(31) => data_im_in(2020),
            data_re_out(0) => first_stage_re_out(36),
            data_re_out(1) => first_stage_re_out(100),
            data_re_out(2) => first_stage_re_out(164),
            data_re_out(3) => first_stage_re_out(228),
            data_re_out(4) => first_stage_re_out(292),
            data_re_out(5) => first_stage_re_out(356),
            data_re_out(6) => first_stage_re_out(420),
            data_re_out(7) => first_stage_re_out(484),
            data_re_out(8) => first_stage_re_out(548),
            data_re_out(9) => first_stage_re_out(612),
            data_re_out(10) => first_stage_re_out(676),
            data_re_out(11) => first_stage_re_out(740),
            data_re_out(12) => first_stage_re_out(804),
            data_re_out(13) => first_stage_re_out(868),
            data_re_out(14) => first_stage_re_out(932),
            data_re_out(15) => first_stage_re_out(996),
            data_re_out(16) => first_stage_re_out(1060),
            data_re_out(17) => first_stage_re_out(1124),
            data_re_out(18) => first_stage_re_out(1188),
            data_re_out(19) => first_stage_re_out(1252),
            data_re_out(20) => first_stage_re_out(1316),
            data_re_out(21) => first_stage_re_out(1380),
            data_re_out(22) => first_stage_re_out(1444),
            data_re_out(23) => first_stage_re_out(1508),
            data_re_out(24) => first_stage_re_out(1572),
            data_re_out(25) => first_stage_re_out(1636),
            data_re_out(26) => first_stage_re_out(1700),
            data_re_out(27) => first_stage_re_out(1764),
            data_re_out(28) => first_stage_re_out(1828),
            data_re_out(29) => first_stage_re_out(1892),
            data_re_out(30) => first_stage_re_out(1956),
            data_re_out(31) => first_stage_re_out(2020),
            data_im_out(0) => first_stage_im_out(36),
            data_im_out(1) => first_stage_im_out(100),
            data_im_out(2) => first_stage_im_out(164),
            data_im_out(3) => first_stage_im_out(228),
            data_im_out(4) => first_stage_im_out(292),
            data_im_out(5) => first_stage_im_out(356),
            data_im_out(6) => first_stage_im_out(420),
            data_im_out(7) => first_stage_im_out(484),
            data_im_out(8) => first_stage_im_out(548),
            data_im_out(9) => first_stage_im_out(612),
            data_im_out(10) => first_stage_im_out(676),
            data_im_out(11) => first_stage_im_out(740),
            data_im_out(12) => first_stage_im_out(804),
            data_im_out(13) => first_stage_im_out(868),
            data_im_out(14) => first_stage_im_out(932),
            data_im_out(15) => first_stage_im_out(996),
            data_im_out(16) => first_stage_im_out(1060),
            data_im_out(17) => first_stage_im_out(1124),
            data_im_out(18) => first_stage_im_out(1188),
            data_im_out(19) => first_stage_im_out(1252),
            data_im_out(20) => first_stage_im_out(1316),
            data_im_out(21) => first_stage_im_out(1380),
            data_im_out(22) => first_stage_im_out(1444),
            data_im_out(23) => first_stage_im_out(1508),
            data_im_out(24) => first_stage_im_out(1572),
            data_im_out(25) => first_stage_im_out(1636),
            data_im_out(26) => first_stage_im_out(1700),
            data_im_out(27) => first_stage_im_out(1764),
            data_im_out(28) => first_stage_im_out(1828),
            data_im_out(29) => first_stage_im_out(1892),
            data_im_out(30) => first_stage_im_out(1956),
            data_im_out(31) => first_stage_im_out(2020)
        );

    ULFFT_PT32_37 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(37),
            data_re_in(1) => data_re_in(101),
            data_re_in(2) => data_re_in(165),
            data_re_in(3) => data_re_in(229),
            data_re_in(4) => data_re_in(293),
            data_re_in(5) => data_re_in(357),
            data_re_in(6) => data_re_in(421),
            data_re_in(7) => data_re_in(485),
            data_re_in(8) => data_re_in(549),
            data_re_in(9) => data_re_in(613),
            data_re_in(10) => data_re_in(677),
            data_re_in(11) => data_re_in(741),
            data_re_in(12) => data_re_in(805),
            data_re_in(13) => data_re_in(869),
            data_re_in(14) => data_re_in(933),
            data_re_in(15) => data_re_in(997),
            data_re_in(16) => data_re_in(1061),
            data_re_in(17) => data_re_in(1125),
            data_re_in(18) => data_re_in(1189),
            data_re_in(19) => data_re_in(1253),
            data_re_in(20) => data_re_in(1317),
            data_re_in(21) => data_re_in(1381),
            data_re_in(22) => data_re_in(1445),
            data_re_in(23) => data_re_in(1509),
            data_re_in(24) => data_re_in(1573),
            data_re_in(25) => data_re_in(1637),
            data_re_in(26) => data_re_in(1701),
            data_re_in(27) => data_re_in(1765),
            data_re_in(28) => data_re_in(1829),
            data_re_in(29) => data_re_in(1893),
            data_re_in(30) => data_re_in(1957),
            data_re_in(31) => data_re_in(2021),
            data_im_in(0) => data_im_in(37),
            data_im_in(1) => data_im_in(101),
            data_im_in(2) => data_im_in(165),
            data_im_in(3) => data_im_in(229),
            data_im_in(4) => data_im_in(293),
            data_im_in(5) => data_im_in(357),
            data_im_in(6) => data_im_in(421),
            data_im_in(7) => data_im_in(485),
            data_im_in(8) => data_im_in(549),
            data_im_in(9) => data_im_in(613),
            data_im_in(10) => data_im_in(677),
            data_im_in(11) => data_im_in(741),
            data_im_in(12) => data_im_in(805),
            data_im_in(13) => data_im_in(869),
            data_im_in(14) => data_im_in(933),
            data_im_in(15) => data_im_in(997),
            data_im_in(16) => data_im_in(1061),
            data_im_in(17) => data_im_in(1125),
            data_im_in(18) => data_im_in(1189),
            data_im_in(19) => data_im_in(1253),
            data_im_in(20) => data_im_in(1317),
            data_im_in(21) => data_im_in(1381),
            data_im_in(22) => data_im_in(1445),
            data_im_in(23) => data_im_in(1509),
            data_im_in(24) => data_im_in(1573),
            data_im_in(25) => data_im_in(1637),
            data_im_in(26) => data_im_in(1701),
            data_im_in(27) => data_im_in(1765),
            data_im_in(28) => data_im_in(1829),
            data_im_in(29) => data_im_in(1893),
            data_im_in(30) => data_im_in(1957),
            data_im_in(31) => data_im_in(2021),
            data_re_out(0) => first_stage_re_out(37),
            data_re_out(1) => first_stage_re_out(101),
            data_re_out(2) => first_stage_re_out(165),
            data_re_out(3) => first_stage_re_out(229),
            data_re_out(4) => first_stage_re_out(293),
            data_re_out(5) => first_stage_re_out(357),
            data_re_out(6) => first_stage_re_out(421),
            data_re_out(7) => first_stage_re_out(485),
            data_re_out(8) => first_stage_re_out(549),
            data_re_out(9) => first_stage_re_out(613),
            data_re_out(10) => first_stage_re_out(677),
            data_re_out(11) => first_stage_re_out(741),
            data_re_out(12) => first_stage_re_out(805),
            data_re_out(13) => first_stage_re_out(869),
            data_re_out(14) => first_stage_re_out(933),
            data_re_out(15) => first_stage_re_out(997),
            data_re_out(16) => first_stage_re_out(1061),
            data_re_out(17) => first_stage_re_out(1125),
            data_re_out(18) => first_stage_re_out(1189),
            data_re_out(19) => first_stage_re_out(1253),
            data_re_out(20) => first_stage_re_out(1317),
            data_re_out(21) => first_stage_re_out(1381),
            data_re_out(22) => first_stage_re_out(1445),
            data_re_out(23) => first_stage_re_out(1509),
            data_re_out(24) => first_stage_re_out(1573),
            data_re_out(25) => first_stage_re_out(1637),
            data_re_out(26) => first_stage_re_out(1701),
            data_re_out(27) => first_stage_re_out(1765),
            data_re_out(28) => first_stage_re_out(1829),
            data_re_out(29) => first_stage_re_out(1893),
            data_re_out(30) => first_stage_re_out(1957),
            data_re_out(31) => first_stage_re_out(2021),
            data_im_out(0) => first_stage_im_out(37),
            data_im_out(1) => first_stage_im_out(101),
            data_im_out(2) => first_stage_im_out(165),
            data_im_out(3) => first_stage_im_out(229),
            data_im_out(4) => first_stage_im_out(293),
            data_im_out(5) => first_stage_im_out(357),
            data_im_out(6) => first_stage_im_out(421),
            data_im_out(7) => first_stage_im_out(485),
            data_im_out(8) => first_stage_im_out(549),
            data_im_out(9) => first_stage_im_out(613),
            data_im_out(10) => first_stage_im_out(677),
            data_im_out(11) => first_stage_im_out(741),
            data_im_out(12) => first_stage_im_out(805),
            data_im_out(13) => first_stage_im_out(869),
            data_im_out(14) => first_stage_im_out(933),
            data_im_out(15) => first_stage_im_out(997),
            data_im_out(16) => first_stage_im_out(1061),
            data_im_out(17) => first_stage_im_out(1125),
            data_im_out(18) => first_stage_im_out(1189),
            data_im_out(19) => first_stage_im_out(1253),
            data_im_out(20) => first_stage_im_out(1317),
            data_im_out(21) => first_stage_im_out(1381),
            data_im_out(22) => first_stage_im_out(1445),
            data_im_out(23) => first_stage_im_out(1509),
            data_im_out(24) => first_stage_im_out(1573),
            data_im_out(25) => first_stage_im_out(1637),
            data_im_out(26) => first_stage_im_out(1701),
            data_im_out(27) => first_stage_im_out(1765),
            data_im_out(28) => first_stage_im_out(1829),
            data_im_out(29) => first_stage_im_out(1893),
            data_im_out(30) => first_stage_im_out(1957),
            data_im_out(31) => first_stage_im_out(2021)
        );

    ULFFT_PT32_38 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(38),
            data_re_in(1) => data_re_in(102),
            data_re_in(2) => data_re_in(166),
            data_re_in(3) => data_re_in(230),
            data_re_in(4) => data_re_in(294),
            data_re_in(5) => data_re_in(358),
            data_re_in(6) => data_re_in(422),
            data_re_in(7) => data_re_in(486),
            data_re_in(8) => data_re_in(550),
            data_re_in(9) => data_re_in(614),
            data_re_in(10) => data_re_in(678),
            data_re_in(11) => data_re_in(742),
            data_re_in(12) => data_re_in(806),
            data_re_in(13) => data_re_in(870),
            data_re_in(14) => data_re_in(934),
            data_re_in(15) => data_re_in(998),
            data_re_in(16) => data_re_in(1062),
            data_re_in(17) => data_re_in(1126),
            data_re_in(18) => data_re_in(1190),
            data_re_in(19) => data_re_in(1254),
            data_re_in(20) => data_re_in(1318),
            data_re_in(21) => data_re_in(1382),
            data_re_in(22) => data_re_in(1446),
            data_re_in(23) => data_re_in(1510),
            data_re_in(24) => data_re_in(1574),
            data_re_in(25) => data_re_in(1638),
            data_re_in(26) => data_re_in(1702),
            data_re_in(27) => data_re_in(1766),
            data_re_in(28) => data_re_in(1830),
            data_re_in(29) => data_re_in(1894),
            data_re_in(30) => data_re_in(1958),
            data_re_in(31) => data_re_in(2022),
            data_im_in(0) => data_im_in(38),
            data_im_in(1) => data_im_in(102),
            data_im_in(2) => data_im_in(166),
            data_im_in(3) => data_im_in(230),
            data_im_in(4) => data_im_in(294),
            data_im_in(5) => data_im_in(358),
            data_im_in(6) => data_im_in(422),
            data_im_in(7) => data_im_in(486),
            data_im_in(8) => data_im_in(550),
            data_im_in(9) => data_im_in(614),
            data_im_in(10) => data_im_in(678),
            data_im_in(11) => data_im_in(742),
            data_im_in(12) => data_im_in(806),
            data_im_in(13) => data_im_in(870),
            data_im_in(14) => data_im_in(934),
            data_im_in(15) => data_im_in(998),
            data_im_in(16) => data_im_in(1062),
            data_im_in(17) => data_im_in(1126),
            data_im_in(18) => data_im_in(1190),
            data_im_in(19) => data_im_in(1254),
            data_im_in(20) => data_im_in(1318),
            data_im_in(21) => data_im_in(1382),
            data_im_in(22) => data_im_in(1446),
            data_im_in(23) => data_im_in(1510),
            data_im_in(24) => data_im_in(1574),
            data_im_in(25) => data_im_in(1638),
            data_im_in(26) => data_im_in(1702),
            data_im_in(27) => data_im_in(1766),
            data_im_in(28) => data_im_in(1830),
            data_im_in(29) => data_im_in(1894),
            data_im_in(30) => data_im_in(1958),
            data_im_in(31) => data_im_in(2022),
            data_re_out(0) => first_stage_re_out(38),
            data_re_out(1) => first_stage_re_out(102),
            data_re_out(2) => first_stage_re_out(166),
            data_re_out(3) => first_stage_re_out(230),
            data_re_out(4) => first_stage_re_out(294),
            data_re_out(5) => first_stage_re_out(358),
            data_re_out(6) => first_stage_re_out(422),
            data_re_out(7) => first_stage_re_out(486),
            data_re_out(8) => first_stage_re_out(550),
            data_re_out(9) => first_stage_re_out(614),
            data_re_out(10) => first_stage_re_out(678),
            data_re_out(11) => first_stage_re_out(742),
            data_re_out(12) => first_stage_re_out(806),
            data_re_out(13) => first_stage_re_out(870),
            data_re_out(14) => first_stage_re_out(934),
            data_re_out(15) => first_stage_re_out(998),
            data_re_out(16) => first_stage_re_out(1062),
            data_re_out(17) => first_stage_re_out(1126),
            data_re_out(18) => first_stage_re_out(1190),
            data_re_out(19) => first_stage_re_out(1254),
            data_re_out(20) => first_stage_re_out(1318),
            data_re_out(21) => first_stage_re_out(1382),
            data_re_out(22) => first_stage_re_out(1446),
            data_re_out(23) => first_stage_re_out(1510),
            data_re_out(24) => first_stage_re_out(1574),
            data_re_out(25) => first_stage_re_out(1638),
            data_re_out(26) => first_stage_re_out(1702),
            data_re_out(27) => first_stage_re_out(1766),
            data_re_out(28) => first_stage_re_out(1830),
            data_re_out(29) => first_stage_re_out(1894),
            data_re_out(30) => first_stage_re_out(1958),
            data_re_out(31) => first_stage_re_out(2022),
            data_im_out(0) => first_stage_im_out(38),
            data_im_out(1) => first_stage_im_out(102),
            data_im_out(2) => first_stage_im_out(166),
            data_im_out(3) => first_stage_im_out(230),
            data_im_out(4) => first_stage_im_out(294),
            data_im_out(5) => first_stage_im_out(358),
            data_im_out(6) => first_stage_im_out(422),
            data_im_out(7) => first_stage_im_out(486),
            data_im_out(8) => first_stage_im_out(550),
            data_im_out(9) => first_stage_im_out(614),
            data_im_out(10) => first_stage_im_out(678),
            data_im_out(11) => first_stage_im_out(742),
            data_im_out(12) => first_stage_im_out(806),
            data_im_out(13) => first_stage_im_out(870),
            data_im_out(14) => first_stage_im_out(934),
            data_im_out(15) => first_stage_im_out(998),
            data_im_out(16) => first_stage_im_out(1062),
            data_im_out(17) => first_stage_im_out(1126),
            data_im_out(18) => first_stage_im_out(1190),
            data_im_out(19) => first_stage_im_out(1254),
            data_im_out(20) => first_stage_im_out(1318),
            data_im_out(21) => first_stage_im_out(1382),
            data_im_out(22) => first_stage_im_out(1446),
            data_im_out(23) => first_stage_im_out(1510),
            data_im_out(24) => first_stage_im_out(1574),
            data_im_out(25) => first_stage_im_out(1638),
            data_im_out(26) => first_stage_im_out(1702),
            data_im_out(27) => first_stage_im_out(1766),
            data_im_out(28) => first_stage_im_out(1830),
            data_im_out(29) => first_stage_im_out(1894),
            data_im_out(30) => first_stage_im_out(1958),
            data_im_out(31) => first_stage_im_out(2022)
        );

    ULFFT_PT32_39 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(39),
            data_re_in(1) => data_re_in(103),
            data_re_in(2) => data_re_in(167),
            data_re_in(3) => data_re_in(231),
            data_re_in(4) => data_re_in(295),
            data_re_in(5) => data_re_in(359),
            data_re_in(6) => data_re_in(423),
            data_re_in(7) => data_re_in(487),
            data_re_in(8) => data_re_in(551),
            data_re_in(9) => data_re_in(615),
            data_re_in(10) => data_re_in(679),
            data_re_in(11) => data_re_in(743),
            data_re_in(12) => data_re_in(807),
            data_re_in(13) => data_re_in(871),
            data_re_in(14) => data_re_in(935),
            data_re_in(15) => data_re_in(999),
            data_re_in(16) => data_re_in(1063),
            data_re_in(17) => data_re_in(1127),
            data_re_in(18) => data_re_in(1191),
            data_re_in(19) => data_re_in(1255),
            data_re_in(20) => data_re_in(1319),
            data_re_in(21) => data_re_in(1383),
            data_re_in(22) => data_re_in(1447),
            data_re_in(23) => data_re_in(1511),
            data_re_in(24) => data_re_in(1575),
            data_re_in(25) => data_re_in(1639),
            data_re_in(26) => data_re_in(1703),
            data_re_in(27) => data_re_in(1767),
            data_re_in(28) => data_re_in(1831),
            data_re_in(29) => data_re_in(1895),
            data_re_in(30) => data_re_in(1959),
            data_re_in(31) => data_re_in(2023),
            data_im_in(0) => data_im_in(39),
            data_im_in(1) => data_im_in(103),
            data_im_in(2) => data_im_in(167),
            data_im_in(3) => data_im_in(231),
            data_im_in(4) => data_im_in(295),
            data_im_in(5) => data_im_in(359),
            data_im_in(6) => data_im_in(423),
            data_im_in(7) => data_im_in(487),
            data_im_in(8) => data_im_in(551),
            data_im_in(9) => data_im_in(615),
            data_im_in(10) => data_im_in(679),
            data_im_in(11) => data_im_in(743),
            data_im_in(12) => data_im_in(807),
            data_im_in(13) => data_im_in(871),
            data_im_in(14) => data_im_in(935),
            data_im_in(15) => data_im_in(999),
            data_im_in(16) => data_im_in(1063),
            data_im_in(17) => data_im_in(1127),
            data_im_in(18) => data_im_in(1191),
            data_im_in(19) => data_im_in(1255),
            data_im_in(20) => data_im_in(1319),
            data_im_in(21) => data_im_in(1383),
            data_im_in(22) => data_im_in(1447),
            data_im_in(23) => data_im_in(1511),
            data_im_in(24) => data_im_in(1575),
            data_im_in(25) => data_im_in(1639),
            data_im_in(26) => data_im_in(1703),
            data_im_in(27) => data_im_in(1767),
            data_im_in(28) => data_im_in(1831),
            data_im_in(29) => data_im_in(1895),
            data_im_in(30) => data_im_in(1959),
            data_im_in(31) => data_im_in(2023),
            data_re_out(0) => first_stage_re_out(39),
            data_re_out(1) => first_stage_re_out(103),
            data_re_out(2) => first_stage_re_out(167),
            data_re_out(3) => first_stage_re_out(231),
            data_re_out(4) => first_stage_re_out(295),
            data_re_out(5) => first_stage_re_out(359),
            data_re_out(6) => first_stage_re_out(423),
            data_re_out(7) => first_stage_re_out(487),
            data_re_out(8) => first_stage_re_out(551),
            data_re_out(9) => first_stage_re_out(615),
            data_re_out(10) => first_stage_re_out(679),
            data_re_out(11) => first_stage_re_out(743),
            data_re_out(12) => first_stage_re_out(807),
            data_re_out(13) => first_stage_re_out(871),
            data_re_out(14) => first_stage_re_out(935),
            data_re_out(15) => first_stage_re_out(999),
            data_re_out(16) => first_stage_re_out(1063),
            data_re_out(17) => first_stage_re_out(1127),
            data_re_out(18) => first_stage_re_out(1191),
            data_re_out(19) => first_stage_re_out(1255),
            data_re_out(20) => first_stage_re_out(1319),
            data_re_out(21) => first_stage_re_out(1383),
            data_re_out(22) => first_stage_re_out(1447),
            data_re_out(23) => first_stage_re_out(1511),
            data_re_out(24) => first_stage_re_out(1575),
            data_re_out(25) => first_stage_re_out(1639),
            data_re_out(26) => first_stage_re_out(1703),
            data_re_out(27) => first_stage_re_out(1767),
            data_re_out(28) => first_stage_re_out(1831),
            data_re_out(29) => first_stage_re_out(1895),
            data_re_out(30) => first_stage_re_out(1959),
            data_re_out(31) => first_stage_re_out(2023),
            data_im_out(0) => first_stage_im_out(39),
            data_im_out(1) => first_stage_im_out(103),
            data_im_out(2) => first_stage_im_out(167),
            data_im_out(3) => first_stage_im_out(231),
            data_im_out(4) => first_stage_im_out(295),
            data_im_out(5) => first_stage_im_out(359),
            data_im_out(6) => first_stage_im_out(423),
            data_im_out(7) => first_stage_im_out(487),
            data_im_out(8) => first_stage_im_out(551),
            data_im_out(9) => first_stage_im_out(615),
            data_im_out(10) => first_stage_im_out(679),
            data_im_out(11) => first_stage_im_out(743),
            data_im_out(12) => first_stage_im_out(807),
            data_im_out(13) => first_stage_im_out(871),
            data_im_out(14) => first_stage_im_out(935),
            data_im_out(15) => first_stage_im_out(999),
            data_im_out(16) => first_stage_im_out(1063),
            data_im_out(17) => first_stage_im_out(1127),
            data_im_out(18) => first_stage_im_out(1191),
            data_im_out(19) => first_stage_im_out(1255),
            data_im_out(20) => first_stage_im_out(1319),
            data_im_out(21) => first_stage_im_out(1383),
            data_im_out(22) => first_stage_im_out(1447),
            data_im_out(23) => first_stage_im_out(1511),
            data_im_out(24) => first_stage_im_out(1575),
            data_im_out(25) => first_stage_im_out(1639),
            data_im_out(26) => first_stage_im_out(1703),
            data_im_out(27) => first_stage_im_out(1767),
            data_im_out(28) => first_stage_im_out(1831),
            data_im_out(29) => first_stage_im_out(1895),
            data_im_out(30) => first_stage_im_out(1959),
            data_im_out(31) => first_stage_im_out(2023)
        );

    ULFFT_PT32_40 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(40),
            data_re_in(1) => data_re_in(104),
            data_re_in(2) => data_re_in(168),
            data_re_in(3) => data_re_in(232),
            data_re_in(4) => data_re_in(296),
            data_re_in(5) => data_re_in(360),
            data_re_in(6) => data_re_in(424),
            data_re_in(7) => data_re_in(488),
            data_re_in(8) => data_re_in(552),
            data_re_in(9) => data_re_in(616),
            data_re_in(10) => data_re_in(680),
            data_re_in(11) => data_re_in(744),
            data_re_in(12) => data_re_in(808),
            data_re_in(13) => data_re_in(872),
            data_re_in(14) => data_re_in(936),
            data_re_in(15) => data_re_in(1000),
            data_re_in(16) => data_re_in(1064),
            data_re_in(17) => data_re_in(1128),
            data_re_in(18) => data_re_in(1192),
            data_re_in(19) => data_re_in(1256),
            data_re_in(20) => data_re_in(1320),
            data_re_in(21) => data_re_in(1384),
            data_re_in(22) => data_re_in(1448),
            data_re_in(23) => data_re_in(1512),
            data_re_in(24) => data_re_in(1576),
            data_re_in(25) => data_re_in(1640),
            data_re_in(26) => data_re_in(1704),
            data_re_in(27) => data_re_in(1768),
            data_re_in(28) => data_re_in(1832),
            data_re_in(29) => data_re_in(1896),
            data_re_in(30) => data_re_in(1960),
            data_re_in(31) => data_re_in(2024),
            data_im_in(0) => data_im_in(40),
            data_im_in(1) => data_im_in(104),
            data_im_in(2) => data_im_in(168),
            data_im_in(3) => data_im_in(232),
            data_im_in(4) => data_im_in(296),
            data_im_in(5) => data_im_in(360),
            data_im_in(6) => data_im_in(424),
            data_im_in(7) => data_im_in(488),
            data_im_in(8) => data_im_in(552),
            data_im_in(9) => data_im_in(616),
            data_im_in(10) => data_im_in(680),
            data_im_in(11) => data_im_in(744),
            data_im_in(12) => data_im_in(808),
            data_im_in(13) => data_im_in(872),
            data_im_in(14) => data_im_in(936),
            data_im_in(15) => data_im_in(1000),
            data_im_in(16) => data_im_in(1064),
            data_im_in(17) => data_im_in(1128),
            data_im_in(18) => data_im_in(1192),
            data_im_in(19) => data_im_in(1256),
            data_im_in(20) => data_im_in(1320),
            data_im_in(21) => data_im_in(1384),
            data_im_in(22) => data_im_in(1448),
            data_im_in(23) => data_im_in(1512),
            data_im_in(24) => data_im_in(1576),
            data_im_in(25) => data_im_in(1640),
            data_im_in(26) => data_im_in(1704),
            data_im_in(27) => data_im_in(1768),
            data_im_in(28) => data_im_in(1832),
            data_im_in(29) => data_im_in(1896),
            data_im_in(30) => data_im_in(1960),
            data_im_in(31) => data_im_in(2024),
            data_re_out(0) => first_stage_re_out(40),
            data_re_out(1) => first_stage_re_out(104),
            data_re_out(2) => first_stage_re_out(168),
            data_re_out(3) => first_stage_re_out(232),
            data_re_out(4) => first_stage_re_out(296),
            data_re_out(5) => first_stage_re_out(360),
            data_re_out(6) => first_stage_re_out(424),
            data_re_out(7) => first_stage_re_out(488),
            data_re_out(8) => first_stage_re_out(552),
            data_re_out(9) => first_stage_re_out(616),
            data_re_out(10) => first_stage_re_out(680),
            data_re_out(11) => first_stage_re_out(744),
            data_re_out(12) => first_stage_re_out(808),
            data_re_out(13) => first_stage_re_out(872),
            data_re_out(14) => first_stage_re_out(936),
            data_re_out(15) => first_stage_re_out(1000),
            data_re_out(16) => first_stage_re_out(1064),
            data_re_out(17) => first_stage_re_out(1128),
            data_re_out(18) => first_stage_re_out(1192),
            data_re_out(19) => first_stage_re_out(1256),
            data_re_out(20) => first_stage_re_out(1320),
            data_re_out(21) => first_stage_re_out(1384),
            data_re_out(22) => first_stage_re_out(1448),
            data_re_out(23) => first_stage_re_out(1512),
            data_re_out(24) => first_stage_re_out(1576),
            data_re_out(25) => first_stage_re_out(1640),
            data_re_out(26) => first_stage_re_out(1704),
            data_re_out(27) => first_stage_re_out(1768),
            data_re_out(28) => first_stage_re_out(1832),
            data_re_out(29) => first_stage_re_out(1896),
            data_re_out(30) => first_stage_re_out(1960),
            data_re_out(31) => first_stage_re_out(2024),
            data_im_out(0) => first_stage_im_out(40),
            data_im_out(1) => first_stage_im_out(104),
            data_im_out(2) => first_stage_im_out(168),
            data_im_out(3) => first_stage_im_out(232),
            data_im_out(4) => first_stage_im_out(296),
            data_im_out(5) => first_stage_im_out(360),
            data_im_out(6) => first_stage_im_out(424),
            data_im_out(7) => first_stage_im_out(488),
            data_im_out(8) => first_stage_im_out(552),
            data_im_out(9) => first_stage_im_out(616),
            data_im_out(10) => first_stage_im_out(680),
            data_im_out(11) => first_stage_im_out(744),
            data_im_out(12) => first_stage_im_out(808),
            data_im_out(13) => first_stage_im_out(872),
            data_im_out(14) => first_stage_im_out(936),
            data_im_out(15) => first_stage_im_out(1000),
            data_im_out(16) => first_stage_im_out(1064),
            data_im_out(17) => first_stage_im_out(1128),
            data_im_out(18) => first_stage_im_out(1192),
            data_im_out(19) => first_stage_im_out(1256),
            data_im_out(20) => first_stage_im_out(1320),
            data_im_out(21) => first_stage_im_out(1384),
            data_im_out(22) => first_stage_im_out(1448),
            data_im_out(23) => first_stage_im_out(1512),
            data_im_out(24) => first_stage_im_out(1576),
            data_im_out(25) => first_stage_im_out(1640),
            data_im_out(26) => first_stage_im_out(1704),
            data_im_out(27) => first_stage_im_out(1768),
            data_im_out(28) => first_stage_im_out(1832),
            data_im_out(29) => first_stage_im_out(1896),
            data_im_out(30) => first_stage_im_out(1960),
            data_im_out(31) => first_stage_im_out(2024)
        );

    ULFFT_PT32_41 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(41),
            data_re_in(1) => data_re_in(105),
            data_re_in(2) => data_re_in(169),
            data_re_in(3) => data_re_in(233),
            data_re_in(4) => data_re_in(297),
            data_re_in(5) => data_re_in(361),
            data_re_in(6) => data_re_in(425),
            data_re_in(7) => data_re_in(489),
            data_re_in(8) => data_re_in(553),
            data_re_in(9) => data_re_in(617),
            data_re_in(10) => data_re_in(681),
            data_re_in(11) => data_re_in(745),
            data_re_in(12) => data_re_in(809),
            data_re_in(13) => data_re_in(873),
            data_re_in(14) => data_re_in(937),
            data_re_in(15) => data_re_in(1001),
            data_re_in(16) => data_re_in(1065),
            data_re_in(17) => data_re_in(1129),
            data_re_in(18) => data_re_in(1193),
            data_re_in(19) => data_re_in(1257),
            data_re_in(20) => data_re_in(1321),
            data_re_in(21) => data_re_in(1385),
            data_re_in(22) => data_re_in(1449),
            data_re_in(23) => data_re_in(1513),
            data_re_in(24) => data_re_in(1577),
            data_re_in(25) => data_re_in(1641),
            data_re_in(26) => data_re_in(1705),
            data_re_in(27) => data_re_in(1769),
            data_re_in(28) => data_re_in(1833),
            data_re_in(29) => data_re_in(1897),
            data_re_in(30) => data_re_in(1961),
            data_re_in(31) => data_re_in(2025),
            data_im_in(0) => data_im_in(41),
            data_im_in(1) => data_im_in(105),
            data_im_in(2) => data_im_in(169),
            data_im_in(3) => data_im_in(233),
            data_im_in(4) => data_im_in(297),
            data_im_in(5) => data_im_in(361),
            data_im_in(6) => data_im_in(425),
            data_im_in(7) => data_im_in(489),
            data_im_in(8) => data_im_in(553),
            data_im_in(9) => data_im_in(617),
            data_im_in(10) => data_im_in(681),
            data_im_in(11) => data_im_in(745),
            data_im_in(12) => data_im_in(809),
            data_im_in(13) => data_im_in(873),
            data_im_in(14) => data_im_in(937),
            data_im_in(15) => data_im_in(1001),
            data_im_in(16) => data_im_in(1065),
            data_im_in(17) => data_im_in(1129),
            data_im_in(18) => data_im_in(1193),
            data_im_in(19) => data_im_in(1257),
            data_im_in(20) => data_im_in(1321),
            data_im_in(21) => data_im_in(1385),
            data_im_in(22) => data_im_in(1449),
            data_im_in(23) => data_im_in(1513),
            data_im_in(24) => data_im_in(1577),
            data_im_in(25) => data_im_in(1641),
            data_im_in(26) => data_im_in(1705),
            data_im_in(27) => data_im_in(1769),
            data_im_in(28) => data_im_in(1833),
            data_im_in(29) => data_im_in(1897),
            data_im_in(30) => data_im_in(1961),
            data_im_in(31) => data_im_in(2025),
            data_re_out(0) => first_stage_re_out(41),
            data_re_out(1) => first_stage_re_out(105),
            data_re_out(2) => first_stage_re_out(169),
            data_re_out(3) => first_stage_re_out(233),
            data_re_out(4) => first_stage_re_out(297),
            data_re_out(5) => first_stage_re_out(361),
            data_re_out(6) => first_stage_re_out(425),
            data_re_out(7) => first_stage_re_out(489),
            data_re_out(8) => first_stage_re_out(553),
            data_re_out(9) => first_stage_re_out(617),
            data_re_out(10) => first_stage_re_out(681),
            data_re_out(11) => first_stage_re_out(745),
            data_re_out(12) => first_stage_re_out(809),
            data_re_out(13) => first_stage_re_out(873),
            data_re_out(14) => first_stage_re_out(937),
            data_re_out(15) => first_stage_re_out(1001),
            data_re_out(16) => first_stage_re_out(1065),
            data_re_out(17) => first_stage_re_out(1129),
            data_re_out(18) => first_stage_re_out(1193),
            data_re_out(19) => first_stage_re_out(1257),
            data_re_out(20) => first_stage_re_out(1321),
            data_re_out(21) => first_stage_re_out(1385),
            data_re_out(22) => first_stage_re_out(1449),
            data_re_out(23) => first_stage_re_out(1513),
            data_re_out(24) => first_stage_re_out(1577),
            data_re_out(25) => first_stage_re_out(1641),
            data_re_out(26) => first_stage_re_out(1705),
            data_re_out(27) => first_stage_re_out(1769),
            data_re_out(28) => first_stage_re_out(1833),
            data_re_out(29) => first_stage_re_out(1897),
            data_re_out(30) => first_stage_re_out(1961),
            data_re_out(31) => first_stage_re_out(2025),
            data_im_out(0) => first_stage_im_out(41),
            data_im_out(1) => first_stage_im_out(105),
            data_im_out(2) => first_stage_im_out(169),
            data_im_out(3) => first_stage_im_out(233),
            data_im_out(4) => first_stage_im_out(297),
            data_im_out(5) => first_stage_im_out(361),
            data_im_out(6) => first_stage_im_out(425),
            data_im_out(7) => first_stage_im_out(489),
            data_im_out(8) => first_stage_im_out(553),
            data_im_out(9) => first_stage_im_out(617),
            data_im_out(10) => first_stage_im_out(681),
            data_im_out(11) => first_stage_im_out(745),
            data_im_out(12) => first_stage_im_out(809),
            data_im_out(13) => first_stage_im_out(873),
            data_im_out(14) => first_stage_im_out(937),
            data_im_out(15) => first_stage_im_out(1001),
            data_im_out(16) => first_stage_im_out(1065),
            data_im_out(17) => first_stage_im_out(1129),
            data_im_out(18) => first_stage_im_out(1193),
            data_im_out(19) => first_stage_im_out(1257),
            data_im_out(20) => first_stage_im_out(1321),
            data_im_out(21) => first_stage_im_out(1385),
            data_im_out(22) => first_stage_im_out(1449),
            data_im_out(23) => first_stage_im_out(1513),
            data_im_out(24) => first_stage_im_out(1577),
            data_im_out(25) => first_stage_im_out(1641),
            data_im_out(26) => first_stage_im_out(1705),
            data_im_out(27) => first_stage_im_out(1769),
            data_im_out(28) => first_stage_im_out(1833),
            data_im_out(29) => first_stage_im_out(1897),
            data_im_out(30) => first_stage_im_out(1961),
            data_im_out(31) => first_stage_im_out(2025)
        );

    ULFFT_PT32_42 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(42),
            data_re_in(1) => data_re_in(106),
            data_re_in(2) => data_re_in(170),
            data_re_in(3) => data_re_in(234),
            data_re_in(4) => data_re_in(298),
            data_re_in(5) => data_re_in(362),
            data_re_in(6) => data_re_in(426),
            data_re_in(7) => data_re_in(490),
            data_re_in(8) => data_re_in(554),
            data_re_in(9) => data_re_in(618),
            data_re_in(10) => data_re_in(682),
            data_re_in(11) => data_re_in(746),
            data_re_in(12) => data_re_in(810),
            data_re_in(13) => data_re_in(874),
            data_re_in(14) => data_re_in(938),
            data_re_in(15) => data_re_in(1002),
            data_re_in(16) => data_re_in(1066),
            data_re_in(17) => data_re_in(1130),
            data_re_in(18) => data_re_in(1194),
            data_re_in(19) => data_re_in(1258),
            data_re_in(20) => data_re_in(1322),
            data_re_in(21) => data_re_in(1386),
            data_re_in(22) => data_re_in(1450),
            data_re_in(23) => data_re_in(1514),
            data_re_in(24) => data_re_in(1578),
            data_re_in(25) => data_re_in(1642),
            data_re_in(26) => data_re_in(1706),
            data_re_in(27) => data_re_in(1770),
            data_re_in(28) => data_re_in(1834),
            data_re_in(29) => data_re_in(1898),
            data_re_in(30) => data_re_in(1962),
            data_re_in(31) => data_re_in(2026),
            data_im_in(0) => data_im_in(42),
            data_im_in(1) => data_im_in(106),
            data_im_in(2) => data_im_in(170),
            data_im_in(3) => data_im_in(234),
            data_im_in(4) => data_im_in(298),
            data_im_in(5) => data_im_in(362),
            data_im_in(6) => data_im_in(426),
            data_im_in(7) => data_im_in(490),
            data_im_in(8) => data_im_in(554),
            data_im_in(9) => data_im_in(618),
            data_im_in(10) => data_im_in(682),
            data_im_in(11) => data_im_in(746),
            data_im_in(12) => data_im_in(810),
            data_im_in(13) => data_im_in(874),
            data_im_in(14) => data_im_in(938),
            data_im_in(15) => data_im_in(1002),
            data_im_in(16) => data_im_in(1066),
            data_im_in(17) => data_im_in(1130),
            data_im_in(18) => data_im_in(1194),
            data_im_in(19) => data_im_in(1258),
            data_im_in(20) => data_im_in(1322),
            data_im_in(21) => data_im_in(1386),
            data_im_in(22) => data_im_in(1450),
            data_im_in(23) => data_im_in(1514),
            data_im_in(24) => data_im_in(1578),
            data_im_in(25) => data_im_in(1642),
            data_im_in(26) => data_im_in(1706),
            data_im_in(27) => data_im_in(1770),
            data_im_in(28) => data_im_in(1834),
            data_im_in(29) => data_im_in(1898),
            data_im_in(30) => data_im_in(1962),
            data_im_in(31) => data_im_in(2026),
            data_re_out(0) => first_stage_re_out(42),
            data_re_out(1) => first_stage_re_out(106),
            data_re_out(2) => first_stage_re_out(170),
            data_re_out(3) => first_stage_re_out(234),
            data_re_out(4) => first_stage_re_out(298),
            data_re_out(5) => first_stage_re_out(362),
            data_re_out(6) => first_stage_re_out(426),
            data_re_out(7) => first_stage_re_out(490),
            data_re_out(8) => first_stage_re_out(554),
            data_re_out(9) => first_stage_re_out(618),
            data_re_out(10) => first_stage_re_out(682),
            data_re_out(11) => first_stage_re_out(746),
            data_re_out(12) => first_stage_re_out(810),
            data_re_out(13) => first_stage_re_out(874),
            data_re_out(14) => first_stage_re_out(938),
            data_re_out(15) => first_stage_re_out(1002),
            data_re_out(16) => first_stage_re_out(1066),
            data_re_out(17) => first_stage_re_out(1130),
            data_re_out(18) => first_stage_re_out(1194),
            data_re_out(19) => first_stage_re_out(1258),
            data_re_out(20) => first_stage_re_out(1322),
            data_re_out(21) => first_stage_re_out(1386),
            data_re_out(22) => first_stage_re_out(1450),
            data_re_out(23) => first_stage_re_out(1514),
            data_re_out(24) => first_stage_re_out(1578),
            data_re_out(25) => first_stage_re_out(1642),
            data_re_out(26) => first_stage_re_out(1706),
            data_re_out(27) => first_stage_re_out(1770),
            data_re_out(28) => first_stage_re_out(1834),
            data_re_out(29) => first_stage_re_out(1898),
            data_re_out(30) => first_stage_re_out(1962),
            data_re_out(31) => first_stage_re_out(2026),
            data_im_out(0) => first_stage_im_out(42),
            data_im_out(1) => first_stage_im_out(106),
            data_im_out(2) => first_stage_im_out(170),
            data_im_out(3) => first_stage_im_out(234),
            data_im_out(4) => first_stage_im_out(298),
            data_im_out(5) => first_stage_im_out(362),
            data_im_out(6) => first_stage_im_out(426),
            data_im_out(7) => first_stage_im_out(490),
            data_im_out(8) => first_stage_im_out(554),
            data_im_out(9) => first_stage_im_out(618),
            data_im_out(10) => first_stage_im_out(682),
            data_im_out(11) => first_stage_im_out(746),
            data_im_out(12) => first_stage_im_out(810),
            data_im_out(13) => first_stage_im_out(874),
            data_im_out(14) => first_stage_im_out(938),
            data_im_out(15) => first_stage_im_out(1002),
            data_im_out(16) => first_stage_im_out(1066),
            data_im_out(17) => first_stage_im_out(1130),
            data_im_out(18) => first_stage_im_out(1194),
            data_im_out(19) => first_stage_im_out(1258),
            data_im_out(20) => first_stage_im_out(1322),
            data_im_out(21) => first_stage_im_out(1386),
            data_im_out(22) => first_stage_im_out(1450),
            data_im_out(23) => first_stage_im_out(1514),
            data_im_out(24) => first_stage_im_out(1578),
            data_im_out(25) => first_stage_im_out(1642),
            data_im_out(26) => first_stage_im_out(1706),
            data_im_out(27) => first_stage_im_out(1770),
            data_im_out(28) => first_stage_im_out(1834),
            data_im_out(29) => first_stage_im_out(1898),
            data_im_out(30) => first_stage_im_out(1962),
            data_im_out(31) => first_stage_im_out(2026)
        );

    ULFFT_PT32_43 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(43),
            data_re_in(1) => data_re_in(107),
            data_re_in(2) => data_re_in(171),
            data_re_in(3) => data_re_in(235),
            data_re_in(4) => data_re_in(299),
            data_re_in(5) => data_re_in(363),
            data_re_in(6) => data_re_in(427),
            data_re_in(7) => data_re_in(491),
            data_re_in(8) => data_re_in(555),
            data_re_in(9) => data_re_in(619),
            data_re_in(10) => data_re_in(683),
            data_re_in(11) => data_re_in(747),
            data_re_in(12) => data_re_in(811),
            data_re_in(13) => data_re_in(875),
            data_re_in(14) => data_re_in(939),
            data_re_in(15) => data_re_in(1003),
            data_re_in(16) => data_re_in(1067),
            data_re_in(17) => data_re_in(1131),
            data_re_in(18) => data_re_in(1195),
            data_re_in(19) => data_re_in(1259),
            data_re_in(20) => data_re_in(1323),
            data_re_in(21) => data_re_in(1387),
            data_re_in(22) => data_re_in(1451),
            data_re_in(23) => data_re_in(1515),
            data_re_in(24) => data_re_in(1579),
            data_re_in(25) => data_re_in(1643),
            data_re_in(26) => data_re_in(1707),
            data_re_in(27) => data_re_in(1771),
            data_re_in(28) => data_re_in(1835),
            data_re_in(29) => data_re_in(1899),
            data_re_in(30) => data_re_in(1963),
            data_re_in(31) => data_re_in(2027),
            data_im_in(0) => data_im_in(43),
            data_im_in(1) => data_im_in(107),
            data_im_in(2) => data_im_in(171),
            data_im_in(3) => data_im_in(235),
            data_im_in(4) => data_im_in(299),
            data_im_in(5) => data_im_in(363),
            data_im_in(6) => data_im_in(427),
            data_im_in(7) => data_im_in(491),
            data_im_in(8) => data_im_in(555),
            data_im_in(9) => data_im_in(619),
            data_im_in(10) => data_im_in(683),
            data_im_in(11) => data_im_in(747),
            data_im_in(12) => data_im_in(811),
            data_im_in(13) => data_im_in(875),
            data_im_in(14) => data_im_in(939),
            data_im_in(15) => data_im_in(1003),
            data_im_in(16) => data_im_in(1067),
            data_im_in(17) => data_im_in(1131),
            data_im_in(18) => data_im_in(1195),
            data_im_in(19) => data_im_in(1259),
            data_im_in(20) => data_im_in(1323),
            data_im_in(21) => data_im_in(1387),
            data_im_in(22) => data_im_in(1451),
            data_im_in(23) => data_im_in(1515),
            data_im_in(24) => data_im_in(1579),
            data_im_in(25) => data_im_in(1643),
            data_im_in(26) => data_im_in(1707),
            data_im_in(27) => data_im_in(1771),
            data_im_in(28) => data_im_in(1835),
            data_im_in(29) => data_im_in(1899),
            data_im_in(30) => data_im_in(1963),
            data_im_in(31) => data_im_in(2027),
            data_re_out(0) => first_stage_re_out(43),
            data_re_out(1) => first_stage_re_out(107),
            data_re_out(2) => first_stage_re_out(171),
            data_re_out(3) => first_stage_re_out(235),
            data_re_out(4) => first_stage_re_out(299),
            data_re_out(5) => first_stage_re_out(363),
            data_re_out(6) => first_stage_re_out(427),
            data_re_out(7) => first_stage_re_out(491),
            data_re_out(8) => first_stage_re_out(555),
            data_re_out(9) => first_stage_re_out(619),
            data_re_out(10) => first_stage_re_out(683),
            data_re_out(11) => first_stage_re_out(747),
            data_re_out(12) => first_stage_re_out(811),
            data_re_out(13) => first_stage_re_out(875),
            data_re_out(14) => first_stage_re_out(939),
            data_re_out(15) => first_stage_re_out(1003),
            data_re_out(16) => first_stage_re_out(1067),
            data_re_out(17) => first_stage_re_out(1131),
            data_re_out(18) => first_stage_re_out(1195),
            data_re_out(19) => first_stage_re_out(1259),
            data_re_out(20) => first_stage_re_out(1323),
            data_re_out(21) => first_stage_re_out(1387),
            data_re_out(22) => first_stage_re_out(1451),
            data_re_out(23) => first_stage_re_out(1515),
            data_re_out(24) => first_stage_re_out(1579),
            data_re_out(25) => first_stage_re_out(1643),
            data_re_out(26) => first_stage_re_out(1707),
            data_re_out(27) => first_stage_re_out(1771),
            data_re_out(28) => first_stage_re_out(1835),
            data_re_out(29) => first_stage_re_out(1899),
            data_re_out(30) => first_stage_re_out(1963),
            data_re_out(31) => first_stage_re_out(2027),
            data_im_out(0) => first_stage_im_out(43),
            data_im_out(1) => first_stage_im_out(107),
            data_im_out(2) => first_stage_im_out(171),
            data_im_out(3) => first_stage_im_out(235),
            data_im_out(4) => first_stage_im_out(299),
            data_im_out(5) => first_stage_im_out(363),
            data_im_out(6) => first_stage_im_out(427),
            data_im_out(7) => first_stage_im_out(491),
            data_im_out(8) => first_stage_im_out(555),
            data_im_out(9) => first_stage_im_out(619),
            data_im_out(10) => first_stage_im_out(683),
            data_im_out(11) => first_stage_im_out(747),
            data_im_out(12) => first_stage_im_out(811),
            data_im_out(13) => first_stage_im_out(875),
            data_im_out(14) => first_stage_im_out(939),
            data_im_out(15) => first_stage_im_out(1003),
            data_im_out(16) => first_stage_im_out(1067),
            data_im_out(17) => first_stage_im_out(1131),
            data_im_out(18) => first_stage_im_out(1195),
            data_im_out(19) => first_stage_im_out(1259),
            data_im_out(20) => first_stage_im_out(1323),
            data_im_out(21) => first_stage_im_out(1387),
            data_im_out(22) => first_stage_im_out(1451),
            data_im_out(23) => first_stage_im_out(1515),
            data_im_out(24) => first_stage_im_out(1579),
            data_im_out(25) => first_stage_im_out(1643),
            data_im_out(26) => first_stage_im_out(1707),
            data_im_out(27) => first_stage_im_out(1771),
            data_im_out(28) => first_stage_im_out(1835),
            data_im_out(29) => first_stage_im_out(1899),
            data_im_out(30) => first_stage_im_out(1963),
            data_im_out(31) => first_stage_im_out(2027)
        );

    ULFFT_PT32_44 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(44),
            data_re_in(1) => data_re_in(108),
            data_re_in(2) => data_re_in(172),
            data_re_in(3) => data_re_in(236),
            data_re_in(4) => data_re_in(300),
            data_re_in(5) => data_re_in(364),
            data_re_in(6) => data_re_in(428),
            data_re_in(7) => data_re_in(492),
            data_re_in(8) => data_re_in(556),
            data_re_in(9) => data_re_in(620),
            data_re_in(10) => data_re_in(684),
            data_re_in(11) => data_re_in(748),
            data_re_in(12) => data_re_in(812),
            data_re_in(13) => data_re_in(876),
            data_re_in(14) => data_re_in(940),
            data_re_in(15) => data_re_in(1004),
            data_re_in(16) => data_re_in(1068),
            data_re_in(17) => data_re_in(1132),
            data_re_in(18) => data_re_in(1196),
            data_re_in(19) => data_re_in(1260),
            data_re_in(20) => data_re_in(1324),
            data_re_in(21) => data_re_in(1388),
            data_re_in(22) => data_re_in(1452),
            data_re_in(23) => data_re_in(1516),
            data_re_in(24) => data_re_in(1580),
            data_re_in(25) => data_re_in(1644),
            data_re_in(26) => data_re_in(1708),
            data_re_in(27) => data_re_in(1772),
            data_re_in(28) => data_re_in(1836),
            data_re_in(29) => data_re_in(1900),
            data_re_in(30) => data_re_in(1964),
            data_re_in(31) => data_re_in(2028),
            data_im_in(0) => data_im_in(44),
            data_im_in(1) => data_im_in(108),
            data_im_in(2) => data_im_in(172),
            data_im_in(3) => data_im_in(236),
            data_im_in(4) => data_im_in(300),
            data_im_in(5) => data_im_in(364),
            data_im_in(6) => data_im_in(428),
            data_im_in(7) => data_im_in(492),
            data_im_in(8) => data_im_in(556),
            data_im_in(9) => data_im_in(620),
            data_im_in(10) => data_im_in(684),
            data_im_in(11) => data_im_in(748),
            data_im_in(12) => data_im_in(812),
            data_im_in(13) => data_im_in(876),
            data_im_in(14) => data_im_in(940),
            data_im_in(15) => data_im_in(1004),
            data_im_in(16) => data_im_in(1068),
            data_im_in(17) => data_im_in(1132),
            data_im_in(18) => data_im_in(1196),
            data_im_in(19) => data_im_in(1260),
            data_im_in(20) => data_im_in(1324),
            data_im_in(21) => data_im_in(1388),
            data_im_in(22) => data_im_in(1452),
            data_im_in(23) => data_im_in(1516),
            data_im_in(24) => data_im_in(1580),
            data_im_in(25) => data_im_in(1644),
            data_im_in(26) => data_im_in(1708),
            data_im_in(27) => data_im_in(1772),
            data_im_in(28) => data_im_in(1836),
            data_im_in(29) => data_im_in(1900),
            data_im_in(30) => data_im_in(1964),
            data_im_in(31) => data_im_in(2028),
            data_re_out(0) => first_stage_re_out(44),
            data_re_out(1) => first_stage_re_out(108),
            data_re_out(2) => first_stage_re_out(172),
            data_re_out(3) => first_stage_re_out(236),
            data_re_out(4) => first_stage_re_out(300),
            data_re_out(5) => first_stage_re_out(364),
            data_re_out(6) => first_stage_re_out(428),
            data_re_out(7) => first_stage_re_out(492),
            data_re_out(8) => first_stage_re_out(556),
            data_re_out(9) => first_stage_re_out(620),
            data_re_out(10) => first_stage_re_out(684),
            data_re_out(11) => first_stage_re_out(748),
            data_re_out(12) => first_stage_re_out(812),
            data_re_out(13) => first_stage_re_out(876),
            data_re_out(14) => first_stage_re_out(940),
            data_re_out(15) => first_stage_re_out(1004),
            data_re_out(16) => first_stage_re_out(1068),
            data_re_out(17) => first_stage_re_out(1132),
            data_re_out(18) => first_stage_re_out(1196),
            data_re_out(19) => first_stage_re_out(1260),
            data_re_out(20) => first_stage_re_out(1324),
            data_re_out(21) => first_stage_re_out(1388),
            data_re_out(22) => first_stage_re_out(1452),
            data_re_out(23) => first_stage_re_out(1516),
            data_re_out(24) => first_stage_re_out(1580),
            data_re_out(25) => first_stage_re_out(1644),
            data_re_out(26) => first_stage_re_out(1708),
            data_re_out(27) => first_stage_re_out(1772),
            data_re_out(28) => first_stage_re_out(1836),
            data_re_out(29) => first_stage_re_out(1900),
            data_re_out(30) => first_stage_re_out(1964),
            data_re_out(31) => first_stage_re_out(2028),
            data_im_out(0) => first_stage_im_out(44),
            data_im_out(1) => first_stage_im_out(108),
            data_im_out(2) => first_stage_im_out(172),
            data_im_out(3) => first_stage_im_out(236),
            data_im_out(4) => first_stage_im_out(300),
            data_im_out(5) => first_stage_im_out(364),
            data_im_out(6) => first_stage_im_out(428),
            data_im_out(7) => first_stage_im_out(492),
            data_im_out(8) => first_stage_im_out(556),
            data_im_out(9) => first_stage_im_out(620),
            data_im_out(10) => first_stage_im_out(684),
            data_im_out(11) => first_stage_im_out(748),
            data_im_out(12) => first_stage_im_out(812),
            data_im_out(13) => first_stage_im_out(876),
            data_im_out(14) => first_stage_im_out(940),
            data_im_out(15) => first_stage_im_out(1004),
            data_im_out(16) => first_stage_im_out(1068),
            data_im_out(17) => first_stage_im_out(1132),
            data_im_out(18) => first_stage_im_out(1196),
            data_im_out(19) => first_stage_im_out(1260),
            data_im_out(20) => first_stage_im_out(1324),
            data_im_out(21) => first_stage_im_out(1388),
            data_im_out(22) => first_stage_im_out(1452),
            data_im_out(23) => first_stage_im_out(1516),
            data_im_out(24) => first_stage_im_out(1580),
            data_im_out(25) => first_stage_im_out(1644),
            data_im_out(26) => first_stage_im_out(1708),
            data_im_out(27) => first_stage_im_out(1772),
            data_im_out(28) => first_stage_im_out(1836),
            data_im_out(29) => first_stage_im_out(1900),
            data_im_out(30) => first_stage_im_out(1964),
            data_im_out(31) => first_stage_im_out(2028)
        );

    ULFFT_PT32_45 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(45),
            data_re_in(1) => data_re_in(109),
            data_re_in(2) => data_re_in(173),
            data_re_in(3) => data_re_in(237),
            data_re_in(4) => data_re_in(301),
            data_re_in(5) => data_re_in(365),
            data_re_in(6) => data_re_in(429),
            data_re_in(7) => data_re_in(493),
            data_re_in(8) => data_re_in(557),
            data_re_in(9) => data_re_in(621),
            data_re_in(10) => data_re_in(685),
            data_re_in(11) => data_re_in(749),
            data_re_in(12) => data_re_in(813),
            data_re_in(13) => data_re_in(877),
            data_re_in(14) => data_re_in(941),
            data_re_in(15) => data_re_in(1005),
            data_re_in(16) => data_re_in(1069),
            data_re_in(17) => data_re_in(1133),
            data_re_in(18) => data_re_in(1197),
            data_re_in(19) => data_re_in(1261),
            data_re_in(20) => data_re_in(1325),
            data_re_in(21) => data_re_in(1389),
            data_re_in(22) => data_re_in(1453),
            data_re_in(23) => data_re_in(1517),
            data_re_in(24) => data_re_in(1581),
            data_re_in(25) => data_re_in(1645),
            data_re_in(26) => data_re_in(1709),
            data_re_in(27) => data_re_in(1773),
            data_re_in(28) => data_re_in(1837),
            data_re_in(29) => data_re_in(1901),
            data_re_in(30) => data_re_in(1965),
            data_re_in(31) => data_re_in(2029),
            data_im_in(0) => data_im_in(45),
            data_im_in(1) => data_im_in(109),
            data_im_in(2) => data_im_in(173),
            data_im_in(3) => data_im_in(237),
            data_im_in(4) => data_im_in(301),
            data_im_in(5) => data_im_in(365),
            data_im_in(6) => data_im_in(429),
            data_im_in(7) => data_im_in(493),
            data_im_in(8) => data_im_in(557),
            data_im_in(9) => data_im_in(621),
            data_im_in(10) => data_im_in(685),
            data_im_in(11) => data_im_in(749),
            data_im_in(12) => data_im_in(813),
            data_im_in(13) => data_im_in(877),
            data_im_in(14) => data_im_in(941),
            data_im_in(15) => data_im_in(1005),
            data_im_in(16) => data_im_in(1069),
            data_im_in(17) => data_im_in(1133),
            data_im_in(18) => data_im_in(1197),
            data_im_in(19) => data_im_in(1261),
            data_im_in(20) => data_im_in(1325),
            data_im_in(21) => data_im_in(1389),
            data_im_in(22) => data_im_in(1453),
            data_im_in(23) => data_im_in(1517),
            data_im_in(24) => data_im_in(1581),
            data_im_in(25) => data_im_in(1645),
            data_im_in(26) => data_im_in(1709),
            data_im_in(27) => data_im_in(1773),
            data_im_in(28) => data_im_in(1837),
            data_im_in(29) => data_im_in(1901),
            data_im_in(30) => data_im_in(1965),
            data_im_in(31) => data_im_in(2029),
            data_re_out(0) => first_stage_re_out(45),
            data_re_out(1) => first_stage_re_out(109),
            data_re_out(2) => first_stage_re_out(173),
            data_re_out(3) => first_stage_re_out(237),
            data_re_out(4) => first_stage_re_out(301),
            data_re_out(5) => first_stage_re_out(365),
            data_re_out(6) => first_stage_re_out(429),
            data_re_out(7) => first_stage_re_out(493),
            data_re_out(8) => first_stage_re_out(557),
            data_re_out(9) => first_stage_re_out(621),
            data_re_out(10) => first_stage_re_out(685),
            data_re_out(11) => first_stage_re_out(749),
            data_re_out(12) => first_stage_re_out(813),
            data_re_out(13) => first_stage_re_out(877),
            data_re_out(14) => first_stage_re_out(941),
            data_re_out(15) => first_stage_re_out(1005),
            data_re_out(16) => first_stage_re_out(1069),
            data_re_out(17) => first_stage_re_out(1133),
            data_re_out(18) => first_stage_re_out(1197),
            data_re_out(19) => first_stage_re_out(1261),
            data_re_out(20) => first_stage_re_out(1325),
            data_re_out(21) => first_stage_re_out(1389),
            data_re_out(22) => first_stage_re_out(1453),
            data_re_out(23) => first_stage_re_out(1517),
            data_re_out(24) => first_stage_re_out(1581),
            data_re_out(25) => first_stage_re_out(1645),
            data_re_out(26) => first_stage_re_out(1709),
            data_re_out(27) => first_stage_re_out(1773),
            data_re_out(28) => first_stage_re_out(1837),
            data_re_out(29) => first_stage_re_out(1901),
            data_re_out(30) => first_stage_re_out(1965),
            data_re_out(31) => first_stage_re_out(2029),
            data_im_out(0) => first_stage_im_out(45),
            data_im_out(1) => first_stage_im_out(109),
            data_im_out(2) => first_stage_im_out(173),
            data_im_out(3) => first_stage_im_out(237),
            data_im_out(4) => first_stage_im_out(301),
            data_im_out(5) => first_stage_im_out(365),
            data_im_out(6) => first_stage_im_out(429),
            data_im_out(7) => first_stage_im_out(493),
            data_im_out(8) => first_stage_im_out(557),
            data_im_out(9) => first_stage_im_out(621),
            data_im_out(10) => first_stage_im_out(685),
            data_im_out(11) => first_stage_im_out(749),
            data_im_out(12) => first_stage_im_out(813),
            data_im_out(13) => first_stage_im_out(877),
            data_im_out(14) => first_stage_im_out(941),
            data_im_out(15) => first_stage_im_out(1005),
            data_im_out(16) => first_stage_im_out(1069),
            data_im_out(17) => first_stage_im_out(1133),
            data_im_out(18) => first_stage_im_out(1197),
            data_im_out(19) => first_stage_im_out(1261),
            data_im_out(20) => first_stage_im_out(1325),
            data_im_out(21) => first_stage_im_out(1389),
            data_im_out(22) => first_stage_im_out(1453),
            data_im_out(23) => first_stage_im_out(1517),
            data_im_out(24) => first_stage_im_out(1581),
            data_im_out(25) => first_stage_im_out(1645),
            data_im_out(26) => first_stage_im_out(1709),
            data_im_out(27) => first_stage_im_out(1773),
            data_im_out(28) => first_stage_im_out(1837),
            data_im_out(29) => first_stage_im_out(1901),
            data_im_out(30) => first_stage_im_out(1965),
            data_im_out(31) => first_stage_im_out(2029)
        );

    ULFFT_PT32_46 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(46),
            data_re_in(1) => data_re_in(110),
            data_re_in(2) => data_re_in(174),
            data_re_in(3) => data_re_in(238),
            data_re_in(4) => data_re_in(302),
            data_re_in(5) => data_re_in(366),
            data_re_in(6) => data_re_in(430),
            data_re_in(7) => data_re_in(494),
            data_re_in(8) => data_re_in(558),
            data_re_in(9) => data_re_in(622),
            data_re_in(10) => data_re_in(686),
            data_re_in(11) => data_re_in(750),
            data_re_in(12) => data_re_in(814),
            data_re_in(13) => data_re_in(878),
            data_re_in(14) => data_re_in(942),
            data_re_in(15) => data_re_in(1006),
            data_re_in(16) => data_re_in(1070),
            data_re_in(17) => data_re_in(1134),
            data_re_in(18) => data_re_in(1198),
            data_re_in(19) => data_re_in(1262),
            data_re_in(20) => data_re_in(1326),
            data_re_in(21) => data_re_in(1390),
            data_re_in(22) => data_re_in(1454),
            data_re_in(23) => data_re_in(1518),
            data_re_in(24) => data_re_in(1582),
            data_re_in(25) => data_re_in(1646),
            data_re_in(26) => data_re_in(1710),
            data_re_in(27) => data_re_in(1774),
            data_re_in(28) => data_re_in(1838),
            data_re_in(29) => data_re_in(1902),
            data_re_in(30) => data_re_in(1966),
            data_re_in(31) => data_re_in(2030),
            data_im_in(0) => data_im_in(46),
            data_im_in(1) => data_im_in(110),
            data_im_in(2) => data_im_in(174),
            data_im_in(3) => data_im_in(238),
            data_im_in(4) => data_im_in(302),
            data_im_in(5) => data_im_in(366),
            data_im_in(6) => data_im_in(430),
            data_im_in(7) => data_im_in(494),
            data_im_in(8) => data_im_in(558),
            data_im_in(9) => data_im_in(622),
            data_im_in(10) => data_im_in(686),
            data_im_in(11) => data_im_in(750),
            data_im_in(12) => data_im_in(814),
            data_im_in(13) => data_im_in(878),
            data_im_in(14) => data_im_in(942),
            data_im_in(15) => data_im_in(1006),
            data_im_in(16) => data_im_in(1070),
            data_im_in(17) => data_im_in(1134),
            data_im_in(18) => data_im_in(1198),
            data_im_in(19) => data_im_in(1262),
            data_im_in(20) => data_im_in(1326),
            data_im_in(21) => data_im_in(1390),
            data_im_in(22) => data_im_in(1454),
            data_im_in(23) => data_im_in(1518),
            data_im_in(24) => data_im_in(1582),
            data_im_in(25) => data_im_in(1646),
            data_im_in(26) => data_im_in(1710),
            data_im_in(27) => data_im_in(1774),
            data_im_in(28) => data_im_in(1838),
            data_im_in(29) => data_im_in(1902),
            data_im_in(30) => data_im_in(1966),
            data_im_in(31) => data_im_in(2030),
            data_re_out(0) => first_stage_re_out(46),
            data_re_out(1) => first_stage_re_out(110),
            data_re_out(2) => first_stage_re_out(174),
            data_re_out(3) => first_stage_re_out(238),
            data_re_out(4) => first_stage_re_out(302),
            data_re_out(5) => first_stage_re_out(366),
            data_re_out(6) => first_stage_re_out(430),
            data_re_out(7) => first_stage_re_out(494),
            data_re_out(8) => first_stage_re_out(558),
            data_re_out(9) => first_stage_re_out(622),
            data_re_out(10) => first_stage_re_out(686),
            data_re_out(11) => first_stage_re_out(750),
            data_re_out(12) => first_stage_re_out(814),
            data_re_out(13) => first_stage_re_out(878),
            data_re_out(14) => first_stage_re_out(942),
            data_re_out(15) => first_stage_re_out(1006),
            data_re_out(16) => first_stage_re_out(1070),
            data_re_out(17) => first_stage_re_out(1134),
            data_re_out(18) => first_stage_re_out(1198),
            data_re_out(19) => first_stage_re_out(1262),
            data_re_out(20) => first_stage_re_out(1326),
            data_re_out(21) => first_stage_re_out(1390),
            data_re_out(22) => first_stage_re_out(1454),
            data_re_out(23) => first_stage_re_out(1518),
            data_re_out(24) => first_stage_re_out(1582),
            data_re_out(25) => first_stage_re_out(1646),
            data_re_out(26) => first_stage_re_out(1710),
            data_re_out(27) => first_stage_re_out(1774),
            data_re_out(28) => first_stage_re_out(1838),
            data_re_out(29) => first_stage_re_out(1902),
            data_re_out(30) => first_stage_re_out(1966),
            data_re_out(31) => first_stage_re_out(2030),
            data_im_out(0) => first_stage_im_out(46),
            data_im_out(1) => first_stage_im_out(110),
            data_im_out(2) => first_stage_im_out(174),
            data_im_out(3) => first_stage_im_out(238),
            data_im_out(4) => first_stage_im_out(302),
            data_im_out(5) => first_stage_im_out(366),
            data_im_out(6) => first_stage_im_out(430),
            data_im_out(7) => first_stage_im_out(494),
            data_im_out(8) => first_stage_im_out(558),
            data_im_out(9) => first_stage_im_out(622),
            data_im_out(10) => first_stage_im_out(686),
            data_im_out(11) => first_stage_im_out(750),
            data_im_out(12) => first_stage_im_out(814),
            data_im_out(13) => first_stage_im_out(878),
            data_im_out(14) => first_stage_im_out(942),
            data_im_out(15) => first_stage_im_out(1006),
            data_im_out(16) => first_stage_im_out(1070),
            data_im_out(17) => first_stage_im_out(1134),
            data_im_out(18) => first_stage_im_out(1198),
            data_im_out(19) => first_stage_im_out(1262),
            data_im_out(20) => first_stage_im_out(1326),
            data_im_out(21) => first_stage_im_out(1390),
            data_im_out(22) => first_stage_im_out(1454),
            data_im_out(23) => first_stage_im_out(1518),
            data_im_out(24) => first_stage_im_out(1582),
            data_im_out(25) => first_stage_im_out(1646),
            data_im_out(26) => first_stage_im_out(1710),
            data_im_out(27) => first_stage_im_out(1774),
            data_im_out(28) => first_stage_im_out(1838),
            data_im_out(29) => first_stage_im_out(1902),
            data_im_out(30) => first_stage_im_out(1966),
            data_im_out(31) => first_stage_im_out(2030)
        );

    ULFFT_PT32_47 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(47),
            data_re_in(1) => data_re_in(111),
            data_re_in(2) => data_re_in(175),
            data_re_in(3) => data_re_in(239),
            data_re_in(4) => data_re_in(303),
            data_re_in(5) => data_re_in(367),
            data_re_in(6) => data_re_in(431),
            data_re_in(7) => data_re_in(495),
            data_re_in(8) => data_re_in(559),
            data_re_in(9) => data_re_in(623),
            data_re_in(10) => data_re_in(687),
            data_re_in(11) => data_re_in(751),
            data_re_in(12) => data_re_in(815),
            data_re_in(13) => data_re_in(879),
            data_re_in(14) => data_re_in(943),
            data_re_in(15) => data_re_in(1007),
            data_re_in(16) => data_re_in(1071),
            data_re_in(17) => data_re_in(1135),
            data_re_in(18) => data_re_in(1199),
            data_re_in(19) => data_re_in(1263),
            data_re_in(20) => data_re_in(1327),
            data_re_in(21) => data_re_in(1391),
            data_re_in(22) => data_re_in(1455),
            data_re_in(23) => data_re_in(1519),
            data_re_in(24) => data_re_in(1583),
            data_re_in(25) => data_re_in(1647),
            data_re_in(26) => data_re_in(1711),
            data_re_in(27) => data_re_in(1775),
            data_re_in(28) => data_re_in(1839),
            data_re_in(29) => data_re_in(1903),
            data_re_in(30) => data_re_in(1967),
            data_re_in(31) => data_re_in(2031),
            data_im_in(0) => data_im_in(47),
            data_im_in(1) => data_im_in(111),
            data_im_in(2) => data_im_in(175),
            data_im_in(3) => data_im_in(239),
            data_im_in(4) => data_im_in(303),
            data_im_in(5) => data_im_in(367),
            data_im_in(6) => data_im_in(431),
            data_im_in(7) => data_im_in(495),
            data_im_in(8) => data_im_in(559),
            data_im_in(9) => data_im_in(623),
            data_im_in(10) => data_im_in(687),
            data_im_in(11) => data_im_in(751),
            data_im_in(12) => data_im_in(815),
            data_im_in(13) => data_im_in(879),
            data_im_in(14) => data_im_in(943),
            data_im_in(15) => data_im_in(1007),
            data_im_in(16) => data_im_in(1071),
            data_im_in(17) => data_im_in(1135),
            data_im_in(18) => data_im_in(1199),
            data_im_in(19) => data_im_in(1263),
            data_im_in(20) => data_im_in(1327),
            data_im_in(21) => data_im_in(1391),
            data_im_in(22) => data_im_in(1455),
            data_im_in(23) => data_im_in(1519),
            data_im_in(24) => data_im_in(1583),
            data_im_in(25) => data_im_in(1647),
            data_im_in(26) => data_im_in(1711),
            data_im_in(27) => data_im_in(1775),
            data_im_in(28) => data_im_in(1839),
            data_im_in(29) => data_im_in(1903),
            data_im_in(30) => data_im_in(1967),
            data_im_in(31) => data_im_in(2031),
            data_re_out(0) => first_stage_re_out(47),
            data_re_out(1) => first_stage_re_out(111),
            data_re_out(2) => first_stage_re_out(175),
            data_re_out(3) => first_stage_re_out(239),
            data_re_out(4) => first_stage_re_out(303),
            data_re_out(5) => first_stage_re_out(367),
            data_re_out(6) => first_stage_re_out(431),
            data_re_out(7) => first_stage_re_out(495),
            data_re_out(8) => first_stage_re_out(559),
            data_re_out(9) => first_stage_re_out(623),
            data_re_out(10) => first_stage_re_out(687),
            data_re_out(11) => first_stage_re_out(751),
            data_re_out(12) => first_stage_re_out(815),
            data_re_out(13) => first_stage_re_out(879),
            data_re_out(14) => first_stage_re_out(943),
            data_re_out(15) => first_stage_re_out(1007),
            data_re_out(16) => first_stage_re_out(1071),
            data_re_out(17) => first_stage_re_out(1135),
            data_re_out(18) => first_stage_re_out(1199),
            data_re_out(19) => first_stage_re_out(1263),
            data_re_out(20) => first_stage_re_out(1327),
            data_re_out(21) => first_stage_re_out(1391),
            data_re_out(22) => first_stage_re_out(1455),
            data_re_out(23) => first_stage_re_out(1519),
            data_re_out(24) => first_stage_re_out(1583),
            data_re_out(25) => first_stage_re_out(1647),
            data_re_out(26) => first_stage_re_out(1711),
            data_re_out(27) => first_stage_re_out(1775),
            data_re_out(28) => first_stage_re_out(1839),
            data_re_out(29) => first_stage_re_out(1903),
            data_re_out(30) => first_stage_re_out(1967),
            data_re_out(31) => first_stage_re_out(2031),
            data_im_out(0) => first_stage_im_out(47),
            data_im_out(1) => first_stage_im_out(111),
            data_im_out(2) => first_stage_im_out(175),
            data_im_out(3) => first_stage_im_out(239),
            data_im_out(4) => first_stage_im_out(303),
            data_im_out(5) => first_stage_im_out(367),
            data_im_out(6) => first_stage_im_out(431),
            data_im_out(7) => first_stage_im_out(495),
            data_im_out(8) => first_stage_im_out(559),
            data_im_out(9) => first_stage_im_out(623),
            data_im_out(10) => first_stage_im_out(687),
            data_im_out(11) => first_stage_im_out(751),
            data_im_out(12) => first_stage_im_out(815),
            data_im_out(13) => first_stage_im_out(879),
            data_im_out(14) => first_stage_im_out(943),
            data_im_out(15) => first_stage_im_out(1007),
            data_im_out(16) => first_stage_im_out(1071),
            data_im_out(17) => first_stage_im_out(1135),
            data_im_out(18) => first_stage_im_out(1199),
            data_im_out(19) => first_stage_im_out(1263),
            data_im_out(20) => first_stage_im_out(1327),
            data_im_out(21) => first_stage_im_out(1391),
            data_im_out(22) => first_stage_im_out(1455),
            data_im_out(23) => first_stage_im_out(1519),
            data_im_out(24) => first_stage_im_out(1583),
            data_im_out(25) => first_stage_im_out(1647),
            data_im_out(26) => first_stage_im_out(1711),
            data_im_out(27) => first_stage_im_out(1775),
            data_im_out(28) => first_stage_im_out(1839),
            data_im_out(29) => first_stage_im_out(1903),
            data_im_out(30) => first_stage_im_out(1967),
            data_im_out(31) => first_stage_im_out(2031)
        );

    ULFFT_PT32_48 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(48),
            data_re_in(1) => data_re_in(112),
            data_re_in(2) => data_re_in(176),
            data_re_in(3) => data_re_in(240),
            data_re_in(4) => data_re_in(304),
            data_re_in(5) => data_re_in(368),
            data_re_in(6) => data_re_in(432),
            data_re_in(7) => data_re_in(496),
            data_re_in(8) => data_re_in(560),
            data_re_in(9) => data_re_in(624),
            data_re_in(10) => data_re_in(688),
            data_re_in(11) => data_re_in(752),
            data_re_in(12) => data_re_in(816),
            data_re_in(13) => data_re_in(880),
            data_re_in(14) => data_re_in(944),
            data_re_in(15) => data_re_in(1008),
            data_re_in(16) => data_re_in(1072),
            data_re_in(17) => data_re_in(1136),
            data_re_in(18) => data_re_in(1200),
            data_re_in(19) => data_re_in(1264),
            data_re_in(20) => data_re_in(1328),
            data_re_in(21) => data_re_in(1392),
            data_re_in(22) => data_re_in(1456),
            data_re_in(23) => data_re_in(1520),
            data_re_in(24) => data_re_in(1584),
            data_re_in(25) => data_re_in(1648),
            data_re_in(26) => data_re_in(1712),
            data_re_in(27) => data_re_in(1776),
            data_re_in(28) => data_re_in(1840),
            data_re_in(29) => data_re_in(1904),
            data_re_in(30) => data_re_in(1968),
            data_re_in(31) => data_re_in(2032),
            data_im_in(0) => data_im_in(48),
            data_im_in(1) => data_im_in(112),
            data_im_in(2) => data_im_in(176),
            data_im_in(3) => data_im_in(240),
            data_im_in(4) => data_im_in(304),
            data_im_in(5) => data_im_in(368),
            data_im_in(6) => data_im_in(432),
            data_im_in(7) => data_im_in(496),
            data_im_in(8) => data_im_in(560),
            data_im_in(9) => data_im_in(624),
            data_im_in(10) => data_im_in(688),
            data_im_in(11) => data_im_in(752),
            data_im_in(12) => data_im_in(816),
            data_im_in(13) => data_im_in(880),
            data_im_in(14) => data_im_in(944),
            data_im_in(15) => data_im_in(1008),
            data_im_in(16) => data_im_in(1072),
            data_im_in(17) => data_im_in(1136),
            data_im_in(18) => data_im_in(1200),
            data_im_in(19) => data_im_in(1264),
            data_im_in(20) => data_im_in(1328),
            data_im_in(21) => data_im_in(1392),
            data_im_in(22) => data_im_in(1456),
            data_im_in(23) => data_im_in(1520),
            data_im_in(24) => data_im_in(1584),
            data_im_in(25) => data_im_in(1648),
            data_im_in(26) => data_im_in(1712),
            data_im_in(27) => data_im_in(1776),
            data_im_in(28) => data_im_in(1840),
            data_im_in(29) => data_im_in(1904),
            data_im_in(30) => data_im_in(1968),
            data_im_in(31) => data_im_in(2032),
            data_re_out(0) => first_stage_re_out(48),
            data_re_out(1) => first_stage_re_out(112),
            data_re_out(2) => first_stage_re_out(176),
            data_re_out(3) => first_stage_re_out(240),
            data_re_out(4) => first_stage_re_out(304),
            data_re_out(5) => first_stage_re_out(368),
            data_re_out(6) => first_stage_re_out(432),
            data_re_out(7) => first_stage_re_out(496),
            data_re_out(8) => first_stage_re_out(560),
            data_re_out(9) => first_stage_re_out(624),
            data_re_out(10) => first_stage_re_out(688),
            data_re_out(11) => first_stage_re_out(752),
            data_re_out(12) => first_stage_re_out(816),
            data_re_out(13) => first_stage_re_out(880),
            data_re_out(14) => first_stage_re_out(944),
            data_re_out(15) => first_stage_re_out(1008),
            data_re_out(16) => first_stage_re_out(1072),
            data_re_out(17) => first_stage_re_out(1136),
            data_re_out(18) => first_stage_re_out(1200),
            data_re_out(19) => first_stage_re_out(1264),
            data_re_out(20) => first_stage_re_out(1328),
            data_re_out(21) => first_stage_re_out(1392),
            data_re_out(22) => first_stage_re_out(1456),
            data_re_out(23) => first_stage_re_out(1520),
            data_re_out(24) => first_stage_re_out(1584),
            data_re_out(25) => first_stage_re_out(1648),
            data_re_out(26) => first_stage_re_out(1712),
            data_re_out(27) => first_stage_re_out(1776),
            data_re_out(28) => first_stage_re_out(1840),
            data_re_out(29) => first_stage_re_out(1904),
            data_re_out(30) => first_stage_re_out(1968),
            data_re_out(31) => first_stage_re_out(2032),
            data_im_out(0) => first_stage_im_out(48),
            data_im_out(1) => first_stage_im_out(112),
            data_im_out(2) => first_stage_im_out(176),
            data_im_out(3) => first_stage_im_out(240),
            data_im_out(4) => first_stage_im_out(304),
            data_im_out(5) => first_stage_im_out(368),
            data_im_out(6) => first_stage_im_out(432),
            data_im_out(7) => first_stage_im_out(496),
            data_im_out(8) => first_stage_im_out(560),
            data_im_out(9) => first_stage_im_out(624),
            data_im_out(10) => first_stage_im_out(688),
            data_im_out(11) => first_stage_im_out(752),
            data_im_out(12) => first_stage_im_out(816),
            data_im_out(13) => first_stage_im_out(880),
            data_im_out(14) => first_stage_im_out(944),
            data_im_out(15) => first_stage_im_out(1008),
            data_im_out(16) => first_stage_im_out(1072),
            data_im_out(17) => first_stage_im_out(1136),
            data_im_out(18) => first_stage_im_out(1200),
            data_im_out(19) => first_stage_im_out(1264),
            data_im_out(20) => first_stage_im_out(1328),
            data_im_out(21) => first_stage_im_out(1392),
            data_im_out(22) => first_stage_im_out(1456),
            data_im_out(23) => first_stage_im_out(1520),
            data_im_out(24) => first_stage_im_out(1584),
            data_im_out(25) => first_stage_im_out(1648),
            data_im_out(26) => first_stage_im_out(1712),
            data_im_out(27) => first_stage_im_out(1776),
            data_im_out(28) => first_stage_im_out(1840),
            data_im_out(29) => first_stage_im_out(1904),
            data_im_out(30) => first_stage_im_out(1968),
            data_im_out(31) => first_stage_im_out(2032)
        );

    ULFFT_PT32_49 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(49),
            data_re_in(1) => data_re_in(113),
            data_re_in(2) => data_re_in(177),
            data_re_in(3) => data_re_in(241),
            data_re_in(4) => data_re_in(305),
            data_re_in(5) => data_re_in(369),
            data_re_in(6) => data_re_in(433),
            data_re_in(7) => data_re_in(497),
            data_re_in(8) => data_re_in(561),
            data_re_in(9) => data_re_in(625),
            data_re_in(10) => data_re_in(689),
            data_re_in(11) => data_re_in(753),
            data_re_in(12) => data_re_in(817),
            data_re_in(13) => data_re_in(881),
            data_re_in(14) => data_re_in(945),
            data_re_in(15) => data_re_in(1009),
            data_re_in(16) => data_re_in(1073),
            data_re_in(17) => data_re_in(1137),
            data_re_in(18) => data_re_in(1201),
            data_re_in(19) => data_re_in(1265),
            data_re_in(20) => data_re_in(1329),
            data_re_in(21) => data_re_in(1393),
            data_re_in(22) => data_re_in(1457),
            data_re_in(23) => data_re_in(1521),
            data_re_in(24) => data_re_in(1585),
            data_re_in(25) => data_re_in(1649),
            data_re_in(26) => data_re_in(1713),
            data_re_in(27) => data_re_in(1777),
            data_re_in(28) => data_re_in(1841),
            data_re_in(29) => data_re_in(1905),
            data_re_in(30) => data_re_in(1969),
            data_re_in(31) => data_re_in(2033),
            data_im_in(0) => data_im_in(49),
            data_im_in(1) => data_im_in(113),
            data_im_in(2) => data_im_in(177),
            data_im_in(3) => data_im_in(241),
            data_im_in(4) => data_im_in(305),
            data_im_in(5) => data_im_in(369),
            data_im_in(6) => data_im_in(433),
            data_im_in(7) => data_im_in(497),
            data_im_in(8) => data_im_in(561),
            data_im_in(9) => data_im_in(625),
            data_im_in(10) => data_im_in(689),
            data_im_in(11) => data_im_in(753),
            data_im_in(12) => data_im_in(817),
            data_im_in(13) => data_im_in(881),
            data_im_in(14) => data_im_in(945),
            data_im_in(15) => data_im_in(1009),
            data_im_in(16) => data_im_in(1073),
            data_im_in(17) => data_im_in(1137),
            data_im_in(18) => data_im_in(1201),
            data_im_in(19) => data_im_in(1265),
            data_im_in(20) => data_im_in(1329),
            data_im_in(21) => data_im_in(1393),
            data_im_in(22) => data_im_in(1457),
            data_im_in(23) => data_im_in(1521),
            data_im_in(24) => data_im_in(1585),
            data_im_in(25) => data_im_in(1649),
            data_im_in(26) => data_im_in(1713),
            data_im_in(27) => data_im_in(1777),
            data_im_in(28) => data_im_in(1841),
            data_im_in(29) => data_im_in(1905),
            data_im_in(30) => data_im_in(1969),
            data_im_in(31) => data_im_in(2033),
            data_re_out(0) => first_stage_re_out(49),
            data_re_out(1) => first_stage_re_out(113),
            data_re_out(2) => first_stage_re_out(177),
            data_re_out(3) => first_stage_re_out(241),
            data_re_out(4) => first_stage_re_out(305),
            data_re_out(5) => first_stage_re_out(369),
            data_re_out(6) => first_stage_re_out(433),
            data_re_out(7) => first_stage_re_out(497),
            data_re_out(8) => first_stage_re_out(561),
            data_re_out(9) => first_stage_re_out(625),
            data_re_out(10) => first_stage_re_out(689),
            data_re_out(11) => first_stage_re_out(753),
            data_re_out(12) => first_stage_re_out(817),
            data_re_out(13) => first_stage_re_out(881),
            data_re_out(14) => first_stage_re_out(945),
            data_re_out(15) => first_stage_re_out(1009),
            data_re_out(16) => first_stage_re_out(1073),
            data_re_out(17) => first_stage_re_out(1137),
            data_re_out(18) => first_stage_re_out(1201),
            data_re_out(19) => first_stage_re_out(1265),
            data_re_out(20) => first_stage_re_out(1329),
            data_re_out(21) => first_stage_re_out(1393),
            data_re_out(22) => first_stage_re_out(1457),
            data_re_out(23) => first_stage_re_out(1521),
            data_re_out(24) => first_stage_re_out(1585),
            data_re_out(25) => first_stage_re_out(1649),
            data_re_out(26) => first_stage_re_out(1713),
            data_re_out(27) => first_stage_re_out(1777),
            data_re_out(28) => first_stage_re_out(1841),
            data_re_out(29) => first_stage_re_out(1905),
            data_re_out(30) => first_stage_re_out(1969),
            data_re_out(31) => first_stage_re_out(2033),
            data_im_out(0) => first_stage_im_out(49),
            data_im_out(1) => first_stage_im_out(113),
            data_im_out(2) => first_stage_im_out(177),
            data_im_out(3) => first_stage_im_out(241),
            data_im_out(4) => first_stage_im_out(305),
            data_im_out(5) => first_stage_im_out(369),
            data_im_out(6) => first_stage_im_out(433),
            data_im_out(7) => first_stage_im_out(497),
            data_im_out(8) => first_stage_im_out(561),
            data_im_out(9) => first_stage_im_out(625),
            data_im_out(10) => first_stage_im_out(689),
            data_im_out(11) => first_stage_im_out(753),
            data_im_out(12) => first_stage_im_out(817),
            data_im_out(13) => first_stage_im_out(881),
            data_im_out(14) => first_stage_im_out(945),
            data_im_out(15) => first_stage_im_out(1009),
            data_im_out(16) => first_stage_im_out(1073),
            data_im_out(17) => first_stage_im_out(1137),
            data_im_out(18) => first_stage_im_out(1201),
            data_im_out(19) => first_stage_im_out(1265),
            data_im_out(20) => first_stage_im_out(1329),
            data_im_out(21) => first_stage_im_out(1393),
            data_im_out(22) => first_stage_im_out(1457),
            data_im_out(23) => first_stage_im_out(1521),
            data_im_out(24) => first_stage_im_out(1585),
            data_im_out(25) => first_stage_im_out(1649),
            data_im_out(26) => first_stage_im_out(1713),
            data_im_out(27) => first_stage_im_out(1777),
            data_im_out(28) => first_stage_im_out(1841),
            data_im_out(29) => first_stage_im_out(1905),
            data_im_out(30) => first_stage_im_out(1969),
            data_im_out(31) => first_stage_im_out(2033)
        );

    ULFFT_PT32_50 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(50),
            data_re_in(1) => data_re_in(114),
            data_re_in(2) => data_re_in(178),
            data_re_in(3) => data_re_in(242),
            data_re_in(4) => data_re_in(306),
            data_re_in(5) => data_re_in(370),
            data_re_in(6) => data_re_in(434),
            data_re_in(7) => data_re_in(498),
            data_re_in(8) => data_re_in(562),
            data_re_in(9) => data_re_in(626),
            data_re_in(10) => data_re_in(690),
            data_re_in(11) => data_re_in(754),
            data_re_in(12) => data_re_in(818),
            data_re_in(13) => data_re_in(882),
            data_re_in(14) => data_re_in(946),
            data_re_in(15) => data_re_in(1010),
            data_re_in(16) => data_re_in(1074),
            data_re_in(17) => data_re_in(1138),
            data_re_in(18) => data_re_in(1202),
            data_re_in(19) => data_re_in(1266),
            data_re_in(20) => data_re_in(1330),
            data_re_in(21) => data_re_in(1394),
            data_re_in(22) => data_re_in(1458),
            data_re_in(23) => data_re_in(1522),
            data_re_in(24) => data_re_in(1586),
            data_re_in(25) => data_re_in(1650),
            data_re_in(26) => data_re_in(1714),
            data_re_in(27) => data_re_in(1778),
            data_re_in(28) => data_re_in(1842),
            data_re_in(29) => data_re_in(1906),
            data_re_in(30) => data_re_in(1970),
            data_re_in(31) => data_re_in(2034),
            data_im_in(0) => data_im_in(50),
            data_im_in(1) => data_im_in(114),
            data_im_in(2) => data_im_in(178),
            data_im_in(3) => data_im_in(242),
            data_im_in(4) => data_im_in(306),
            data_im_in(5) => data_im_in(370),
            data_im_in(6) => data_im_in(434),
            data_im_in(7) => data_im_in(498),
            data_im_in(8) => data_im_in(562),
            data_im_in(9) => data_im_in(626),
            data_im_in(10) => data_im_in(690),
            data_im_in(11) => data_im_in(754),
            data_im_in(12) => data_im_in(818),
            data_im_in(13) => data_im_in(882),
            data_im_in(14) => data_im_in(946),
            data_im_in(15) => data_im_in(1010),
            data_im_in(16) => data_im_in(1074),
            data_im_in(17) => data_im_in(1138),
            data_im_in(18) => data_im_in(1202),
            data_im_in(19) => data_im_in(1266),
            data_im_in(20) => data_im_in(1330),
            data_im_in(21) => data_im_in(1394),
            data_im_in(22) => data_im_in(1458),
            data_im_in(23) => data_im_in(1522),
            data_im_in(24) => data_im_in(1586),
            data_im_in(25) => data_im_in(1650),
            data_im_in(26) => data_im_in(1714),
            data_im_in(27) => data_im_in(1778),
            data_im_in(28) => data_im_in(1842),
            data_im_in(29) => data_im_in(1906),
            data_im_in(30) => data_im_in(1970),
            data_im_in(31) => data_im_in(2034),
            data_re_out(0) => first_stage_re_out(50),
            data_re_out(1) => first_stage_re_out(114),
            data_re_out(2) => first_stage_re_out(178),
            data_re_out(3) => first_stage_re_out(242),
            data_re_out(4) => first_stage_re_out(306),
            data_re_out(5) => first_stage_re_out(370),
            data_re_out(6) => first_stage_re_out(434),
            data_re_out(7) => first_stage_re_out(498),
            data_re_out(8) => first_stage_re_out(562),
            data_re_out(9) => first_stage_re_out(626),
            data_re_out(10) => first_stage_re_out(690),
            data_re_out(11) => first_stage_re_out(754),
            data_re_out(12) => first_stage_re_out(818),
            data_re_out(13) => first_stage_re_out(882),
            data_re_out(14) => first_stage_re_out(946),
            data_re_out(15) => first_stage_re_out(1010),
            data_re_out(16) => first_stage_re_out(1074),
            data_re_out(17) => first_stage_re_out(1138),
            data_re_out(18) => first_stage_re_out(1202),
            data_re_out(19) => first_stage_re_out(1266),
            data_re_out(20) => first_stage_re_out(1330),
            data_re_out(21) => first_stage_re_out(1394),
            data_re_out(22) => first_stage_re_out(1458),
            data_re_out(23) => first_stage_re_out(1522),
            data_re_out(24) => first_stage_re_out(1586),
            data_re_out(25) => first_stage_re_out(1650),
            data_re_out(26) => first_stage_re_out(1714),
            data_re_out(27) => first_stage_re_out(1778),
            data_re_out(28) => first_stage_re_out(1842),
            data_re_out(29) => first_stage_re_out(1906),
            data_re_out(30) => first_stage_re_out(1970),
            data_re_out(31) => first_stage_re_out(2034),
            data_im_out(0) => first_stage_im_out(50),
            data_im_out(1) => first_stage_im_out(114),
            data_im_out(2) => first_stage_im_out(178),
            data_im_out(3) => first_stage_im_out(242),
            data_im_out(4) => first_stage_im_out(306),
            data_im_out(5) => first_stage_im_out(370),
            data_im_out(6) => first_stage_im_out(434),
            data_im_out(7) => first_stage_im_out(498),
            data_im_out(8) => first_stage_im_out(562),
            data_im_out(9) => first_stage_im_out(626),
            data_im_out(10) => first_stage_im_out(690),
            data_im_out(11) => first_stage_im_out(754),
            data_im_out(12) => first_stage_im_out(818),
            data_im_out(13) => first_stage_im_out(882),
            data_im_out(14) => first_stage_im_out(946),
            data_im_out(15) => first_stage_im_out(1010),
            data_im_out(16) => first_stage_im_out(1074),
            data_im_out(17) => first_stage_im_out(1138),
            data_im_out(18) => first_stage_im_out(1202),
            data_im_out(19) => first_stage_im_out(1266),
            data_im_out(20) => first_stage_im_out(1330),
            data_im_out(21) => first_stage_im_out(1394),
            data_im_out(22) => first_stage_im_out(1458),
            data_im_out(23) => first_stage_im_out(1522),
            data_im_out(24) => first_stage_im_out(1586),
            data_im_out(25) => first_stage_im_out(1650),
            data_im_out(26) => first_stage_im_out(1714),
            data_im_out(27) => first_stage_im_out(1778),
            data_im_out(28) => first_stage_im_out(1842),
            data_im_out(29) => first_stage_im_out(1906),
            data_im_out(30) => first_stage_im_out(1970),
            data_im_out(31) => first_stage_im_out(2034)
        );

    ULFFT_PT32_51 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(51),
            data_re_in(1) => data_re_in(115),
            data_re_in(2) => data_re_in(179),
            data_re_in(3) => data_re_in(243),
            data_re_in(4) => data_re_in(307),
            data_re_in(5) => data_re_in(371),
            data_re_in(6) => data_re_in(435),
            data_re_in(7) => data_re_in(499),
            data_re_in(8) => data_re_in(563),
            data_re_in(9) => data_re_in(627),
            data_re_in(10) => data_re_in(691),
            data_re_in(11) => data_re_in(755),
            data_re_in(12) => data_re_in(819),
            data_re_in(13) => data_re_in(883),
            data_re_in(14) => data_re_in(947),
            data_re_in(15) => data_re_in(1011),
            data_re_in(16) => data_re_in(1075),
            data_re_in(17) => data_re_in(1139),
            data_re_in(18) => data_re_in(1203),
            data_re_in(19) => data_re_in(1267),
            data_re_in(20) => data_re_in(1331),
            data_re_in(21) => data_re_in(1395),
            data_re_in(22) => data_re_in(1459),
            data_re_in(23) => data_re_in(1523),
            data_re_in(24) => data_re_in(1587),
            data_re_in(25) => data_re_in(1651),
            data_re_in(26) => data_re_in(1715),
            data_re_in(27) => data_re_in(1779),
            data_re_in(28) => data_re_in(1843),
            data_re_in(29) => data_re_in(1907),
            data_re_in(30) => data_re_in(1971),
            data_re_in(31) => data_re_in(2035),
            data_im_in(0) => data_im_in(51),
            data_im_in(1) => data_im_in(115),
            data_im_in(2) => data_im_in(179),
            data_im_in(3) => data_im_in(243),
            data_im_in(4) => data_im_in(307),
            data_im_in(5) => data_im_in(371),
            data_im_in(6) => data_im_in(435),
            data_im_in(7) => data_im_in(499),
            data_im_in(8) => data_im_in(563),
            data_im_in(9) => data_im_in(627),
            data_im_in(10) => data_im_in(691),
            data_im_in(11) => data_im_in(755),
            data_im_in(12) => data_im_in(819),
            data_im_in(13) => data_im_in(883),
            data_im_in(14) => data_im_in(947),
            data_im_in(15) => data_im_in(1011),
            data_im_in(16) => data_im_in(1075),
            data_im_in(17) => data_im_in(1139),
            data_im_in(18) => data_im_in(1203),
            data_im_in(19) => data_im_in(1267),
            data_im_in(20) => data_im_in(1331),
            data_im_in(21) => data_im_in(1395),
            data_im_in(22) => data_im_in(1459),
            data_im_in(23) => data_im_in(1523),
            data_im_in(24) => data_im_in(1587),
            data_im_in(25) => data_im_in(1651),
            data_im_in(26) => data_im_in(1715),
            data_im_in(27) => data_im_in(1779),
            data_im_in(28) => data_im_in(1843),
            data_im_in(29) => data_im_in(1907),
            data_im_in(30) => data_im_in(1971),
            data_im_in(31) => data_im_in(2035),
            data_re_out(0) => first_stage_re_out(51),
            data_re_out(1) => first_stage_re_out(115),
            data_re_out(2) => first_stage_re_out(179),
            data_re_out(3) => first_stage_re_out(243),
            data_re_out(4) => first_stage_re_out(307),
            data_re_out(5) => first_stage_re_out(371),
            data_re_out(6) => first_stage_re_out(435),
            data_re_out(7) => first_stage_re_out(499),
            data_re_out(8) => first_stage_re_out(563),
            data_re_out(9) => first_stage_re_out(627),
            data_re_out(10) => first_stage_re_out(691),
            data_re_out(11) => first_stage_re_out(755),
            data_re_out(12) => first_stage_re_out(819),
            data_re_out(13) => first_stage_re_out(883),
            data_re_out(14) => first_stage_re_out(947),
            data_re_out(15) => first_stage_re_out(1011),
            data_re_out(16) => first_stage_re_out(1075),
            data_re_out(17) => first_stage_re_out(1139),
            data_re_out(18) => first_stage_re_out(1203),
            data_re_out(19) => first_stage_re_out(1267),
            data_re_out(20) => first_stage_re_out(1331),
            data_re_out(21) => first_stage_re_out(1395),
            data_re_out(22) => first_stage_re_out(1459),
            data_re_out(23) => first_stage_re_out(1523),
            data_re_out(24) => first_stage_re_out(1587),
            data_re_out(25) => first_stage_re_out(1651),
            data_re_out(26) => first_stage_re_out(1715),
            data_re_out(27) => first_stage_re_out(1779),
            data_re_out(28) => first_stage_re_out(1843),
            data_re_out(29) => first_stage_re_out(1907),
            data_re_out(30) => first_stage_re_out(1971),
            data_re_out(31) => first_stage_re_out(2035),
            data_im_out(0) => first_stage_im_out(51),
            data_im_out(1) => first_stage_im_out(115),
            data_im_out(2) => first_stage_im_out(179),
            data_im_out(3) => first_stage_im_out(243),
            data_im_out(4) => first_stage_im_out(307),
            data_im_out(5) => first_stage_im_out(371),
            data_im_out(6) => first_stage_im_out(435),
            data_im_out(7) => first_stage_im_out(499),
            data_im_out(8) => first_stage_im_out(563),
            data_im_out(9) => first_stage_im_out(627),
            data_im_out(10) => first_stage_im_out(691),
            data_im_out(11) => first_stage_im_out(755),
            data_im_out(12) => first_stage_im_out(819),
            data_im_out(13) => first_stage_im_out(883),
            data_im_out(14) => first_stage_im_out(947),
            data_im_out(15) => first_stage_im_out(1011),
            data_im_out(16) => first_stage_im_out(1075),
            data_im_out(17) => first_stage_im_out(1139),
            data_im_out(18) => first_stage_im_out(1203),
            data_im_out(19) => first_stage_im_out(1267),
            data_im_out(20) => first_stage_im_out(1331),
            data_im_out(21) => first_stage_im_out(1395),
            data_im_out(22) => first_stage_im_out(1459),
            data_im_out(23) => first_stage_im_out(1523),
            data_im_out(24) => first_stage_im_out(1587),
            data_im_out(25) => first_stage_im_out(1651),
            data_im_out(26) => first_stage_im_out(1715),
            data_im_out(27) => first_stage_im_out(1779),
            data_im_out(28) => first_stage_im_out(1843),
            data_im_out(29) => first_stage_im_out(1907),
            data_im_out(30) => first_stage_im_out(1971),
            data_im_out(31) => first_stage_im_out(2035)
        );

    ULFFT_PT32_52 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(52),
            data_re_in(1) => data_re_in(116),
            data_re_in(2) => data_re_in(180),
            data_re_in(3) => data_re_in(244),
            data_re_in(4) => data_re_in(308),
            data_re_in(5) => data_re_in(372),
            data_re_in(6) => data_re_in(436),
            data_re_in(7) => data_re_in(500),
            data_re_in(8) => data_re_in(564),
            data_re_in(9) => data_re_in(628),
            data_re_in(10) => data_re_in(692),
            data_re_in(11) => data_re_in(756),
            data_re_in(12) => data_re_in(820),
            data_re_in(13) => data_re_in(884),
            data_re_in(14) => data_re_in(948),
            data_re_in(15) => data_re_in(1012),
            data_re_in(16) => data_re_in(1076),
            data_re_in(17) => data_re_in(1140),
            data_re_in(18) => data_re_in(1204),
            data_re_in(19) => data_re_in(1268),
            data_re_in(20) => data_re_in(1332),
            data_re_in(21) => data_re_in(1396),
            data_re_in(22) => data_re_in(1460),
            data_re_in(23) => data_re_in(1524),
            data_re_in(24) => data_re_in(1588),
            data_re_in(25) => data_re_in(1652),
            data_re_in(26) => data_re_in(1716),
            data_re_in(27) => data_re_in(1780),
            data_re_in(28) => data_re_in(1844),
            data_re_in(29) => data_re_in(1908),
            data_re_in(30) => data_re_in(1972),
            data_re_in(31) => data_re_in(2036),
            data_im_in(0) => data_im_in(52),
            data_im_in(1) => data_im_in(116),
            data_im_in(2) => data_im_in(180),
            data_im_in(3) => data_im_in(244),
            data_im_in(4) => data_im_in(308),
            data_im_in(5) => data_im_in(372),
            data_im_in(6) => data_im_in(436),
            data_im_in(7) => data_im_in(500),
            data_im_in(8) => data_im_in(564),
            data_im_in(9) => data_im_in(628),
            data_im_in(10) => data_im_in(692),
            data_im_in(11) => data_im_in(756),
            data_im_in(12) => data_im_in(820),
            data_im_in(13) => data_im_in(884),
            data_im_in(14) => data_im_in(948),
            data_im_in(15) => data_im_in(1012),
            data_im_in(16) => data_im_in(1076),
            data_im_in(17) => data_im_in(1140),
            data_im_in(18) => data_im_in(1204),
            data_im_in(19) => data_im_in(1268),
            data_im_in(20) => data_im_in(1332),
            data_im_in(21) => data_im_in(1396),
            data_im_in(22) => data_im_in(1460),
            data_im_in(23) => data_im_in(1524),
            data_im_in(24) => data_im_in(1588),
            data_im_in(25) => data_im_in(1652),
            data_im_in(26) => data_im_in(1716),
            data_im_in(27) => data_im_in(1780),
            data_im_in(28) => data_im_in(1844),
            data_im_in(29) => data_im_in(1908),
            data_im_in(30) => data_im_in(1972),
            data_im_in(31) => data_im_in(2036),
            data_re_out(0) => first_stage_re_out(52),
            data_re_out(1) => first_stage_re_out(116),
            data_re_out(2) => first_stage_re_out(180),
            data_re_out(3) => first_stage_re_out(244),
            data_re_out(4) => first_stage_re_out(308),
            data_re_out(5) => first_stage_re_out(372),
            data_re_out(6) => first_stage_re_out(436),
            data_re_out(7) => first_stage_re_out(500),
            data_re_out(8) => first_stage_re_out(564),
            data_re_out(9) => first_stage_re_out(628),
            data_re_out(10) => first_stage_re_out(692),
            data_re_out(11) => first_stage_re_out(756),
            data_re_out(12) => first_stage_re_out(820),
            data_re_out(13) => first_stage_re_out(884),
            data_re_out(14) => first_stage_re_out(948),
            data_re_out(15) => first_stage_re_out(1012),
            data_re_out(16) => first_stage_re_out(1076),
            data_re_out(17) => first_stage_re_out(1140),
            data_re_out(18) => first_stage_re_out(1204),
            data_re_out(19) => first_stage_re_out(1268),
            data_re_out(20) => first_stage_re_out(1332),
            data_re_out(21) => first_stage_re_out(1396),
            data_re_out(22) => first_stage_re_out(1460),
            data_re_out(23) => first_stage_re_out(1524),
            data_re_out(24) => first_stage_re_out(1588),
            data_re_out(25) => first_stage_re_out(1652),
            data_re_out(26) => first_stage_re_out(1716),
            data_re_out(27) => first_stage_re_out(1780),
            data_re_out(28) => first_stage_re_out(1844),
            data_re_out(29) => first_stage_re_out(1908),
            data_re_out(30) => first_stage_re_out(1972),
            data_re_out(31) => first_stage_re_out(2036),
            data_im_out(0) => first_stage_im_out(52),
            data_im_out(1) => first_stage_im_out(116),
            data_im_out(2) => first_stage_im_out(180),
            data_im_out(3) => first_stage_im_out(244),
            data_im_out(4) => first_stage_im_out(308),
            data_im_out(5) => first_stage_im_out(372),
            data_im_out(6) => first_stage_im_out(436),
            data_im_out(7) => first_stage_im_out(500),
            data_im_out(8) => first_stage_im_out(564),
            data_im_out(9) => first_stage_im_out(628),
            data_im_out(10) => first_stage_im_out(692),
            data_im_out(11) => first_stage_im_out(756),
            data_im_out(12) => first_stage_im_out(820),
            data_im_out(13) => first_stage_im_out(884),
            data_im_out(14) => first_stage_im_out(948),
            data_im_out(15) => first_stage_im_out(1012),
            data_im_out(16) => first_stage_im_out(1076),
            data_im_out(17) => first_stage_im_out(1140),
            data_im_out(18) => first_stage_im_out(1204),
            data_im_out(19) => first_stage_im_out(1268),
            data_im_out(20) => first_stage_im_out(1332),
            data_im_out(21) => first_stage_im_out(1396),
            data_im_out(22) => first_stage_im_out(1460),
            data_im_out(23) => first_stage_im_out(1524),
            data_im_out(24) => first_stage_im_out(1588),
            data_im_out(25) => first_stage_im_out(1652),
            data_im_out(26) => first_stage_im_out(1716),
            data_im_out(27) => first_stage_im_out(1780),
            data_im_out(28) => first_stage_im_out(1844),
            data_im_out(29) => first_stage_im_out(1908),
            data_im_out(30) => first_stage_im_out(1972),
            data_im_out(31) => first_stage_im_out(2036)
        );

    ULFFT_PT32_53 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(53),
            data_re_in(1) => data_re_in(117),
            data_re_in(2) => data_re_in(181),
            data_re_in(3) => data_re_in(245),
            data_re_in(4) => data_re_in(309),
            data_re_in(5) => data_re_in(373),
            data_re_in(6) => data_re_in(437),
            data_re_in(7) => data_re_in(501),
            data_re_in(8) => data_re_in(565),
            data_re_in(9) => data_re_in(629),
            data_re_in(10) => data_re_in(693),
            data_re_in(11) => data_re_in(757),
            data_re_in(12) => data_re_in(821),
            data_re_in(13) => data_re_in(885),
            data_re_in(14) => data_re_in(949),
            data_re_in(15) => data_re_in(1013),
            data_re_in(16) => data_re_in(1077),
            data_re_in(17) => data_re_in(1141),
            data_re_in(18) => data_re_in(1205),
            data_re_in(19) => data_re_in(1269),
            data_re_in(20) => data_re_in(1333),
            data_re_in(21) => data_re_in(1397),
            data_re_in(22) => data_re_in(1461),
            data_re_in(23) => data_re_in(1525),
            data_re_in(24) => data_re_in(1589),
            data_re_in(25) => data_re_in(1653),
            data_re_in(26) => data_re_in(1717),
            data_re_in(27) => data_re_in(1781),
            data_re_in(28) => data_re_in(1845),
            data_re_in(29) => data_re_in(1909),
            data_re_in(30) => data_re_in(1973),
            data_re_in(31) => data_re_in(2037),
            data_im_in(0) => data_im_in(53),
            data_im_in(1) => data_im_in(117),
            data_im_in(2) => data_im_in(181),
            data_im_in(3) => data_im_in(245),
            data_im_in(4) => data_im_in(309),
            data_im_in(5) => data_im_in(373),
            data_im_in(6) => data_im_in(437),
            data_im_in(7) => data_im_in(501),
            data_im_in(8) => data_im_in(565),
            data_im_in(9) => data_im_in(629),
            data_im_in(10) => data_im_in(693),
            data_im_in(11) => data_im_in(757),
            data_im_in(12) => data_im_in(821),
            data_im_in(13) => data_im_in(885),
            data_im_in(14) => data_im_in(949),
            data_im_in(15) => data_im_in(1013),
            data_im_in(16) => data_im_in(1077),
            data_im_in(17) => data_im_in(1141),
            data_im_in(18) => data_im_in(1205),
            data_im_in(19) => data_im_in(1269),
            data_im_in(20) => data_im_in(1333),
            data_im_in(21) => data_im_in(1397),
            data_im_in(22) => data_im_in(1461),
            data_im_in(23) => data_im_in(1525),
            data_im_in(24) => data_im_in(1589),
            data_im_in(25) => data_im_in(1653),
            data_im_in(26) => data_im_in(1717),
            data_im_in(27) => data_im_in(1781),
            data_im_in(28) => data_im_in(1845),
            data_im_in(29) => data_im_in(1909),
            data_im_in(30) => data_im_in(1973),
            data_im_in(31) => data_im_in(2037),
            data_re_out(0) => first_stage_re_out(53),
            data_re_out(1) => first_stage_re_out(117),
            data_re_out(2) => first_stage_re_out(181),
            data_re_out(3) => first_stage_re_out(245),
            data_re_out(4) => first_stage_re_out(309),
            data_re_out(5) => first_stage_re_out(373),
            data_re_out(6) => first_stage_re_out(437),
            data_re_out(7) => first_stage_re_out(501),
            data_re_out(8) => first_stage_re_out(565),
            data_re_out(9) => first_stage_re_out(629),
            data_re_out(10) => first_stage_re_out(693),
            data_re_out(11) => first_stage_re_out(757),
            data_re_out(12) => first_stage_re_out(821),
            data_re_out(13) => first_stage_re_out(885),
            data_re_out(14) => first_stage_re_out(949),
            data_re_out(15) => first_stage_re_out(1013),
            data_re_out(16) => first_stage_re_out(1077),
            data_re_out(17) => first_stage_re_out(1141),
            data_re_out(18) => first_stage_re_out(1205),
            data_re_out(19) => first_stage_re_out(1269),
            data_re_out(20) => first_stage_re_out(1333),
            data_re_out(21) => first_stage_re_out(1397),
            data_re_out(22) => first_stage_re_out(1461),
            data_re_out(23) => first_stage_re_out(1525),
            data_re_out(24) => first_stage_re_out(1589),
            data_re_out(25) => first_stage_re_out(1653),
            data_re_out(26) => first_stage_re_out(1717),
            data_re_out(27) => first_stage_re_out(1781),
            data_re_out(28) => first_stage_re_out(1845),
            data_re_out(29) => first_stage_re_out(1909),
            data_re_out(30) => first_stage_re_out(1973),
            data_re_out(31) => first_stage_re_out(2037),
            data_im_out(0) => first_stage_im_out(53),
            data_im_out(1) => first_stage_im_out(117),
            data_im_out(2) => first_stage_im_out(181),
            data_im_out(3) => first_stage_im_out(245),
            data_im_out(4) => first_stage_im_out(309),
            data_im_out(5) => first_stage_im_out(373),
            data_im_out(6) => first_stage_im_out(437),
            data_im_out(7) => first_stage_im_out(501),
            data_im_out(8) => first_stage_im_out(565),
            data_im_out(9) => first_stage_im_out(629),
            data_im_out(10) => first_stage_im_out(693),
            data_im_out(11) => first_stage_im_out(757),
            data_im_out(12) => first_stage_im_out(821),
            data_im_out(13) => first_stage_im_out(885),
            data_im_out(14) => first_stage_im_out(949),
            data_im_out(15) => first_stage_im_out(1013),
            data_im_out(16) => first_stage_im_out(1077),
            data_im_out(17) => first_stage_im_out(1141),
            data_im_out(18) => first_stage_im_out(1205),
            data_im_out(19) => first_stage_im_out(1269),
            data_im_out(20) => first_stage_im_out(1333),
            data_im_out(21) => first_stage_im_out(1397),
            data_im_out(22) => first_stage_im_out(1461),
            data_im_out(23) => first_stage_im_out(1525),
            data_im_out(24) => first_stage_im_out(1589),
            data_im_out(25) => first_stage_im_out(1653),
            data_im_out(26) => first_stage_im_out(1717),
            data_im_out(27) => first_stage_im_out(1781),
            data_im_out(28) => first_stage_im_out(1845),
            data_im_out(29) => first_stage_im_out(1909),
            data_im_out(30) => first_stage_im_out(1973),
            data_im_out(31) => first_stage_im_out(2037)
        );

    ULFFT_PT32_54 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(54),
            data_re_in(1) => data_re_in(118),
            data_re_in(2) => data_re_in(182),
            data_re_in(3) => data_re_in(246),
            data_re_in(4) => data_re_in(310),
            data_re_in(5) => data_re_in(374),
            data_re_in(6) => data_re_in(438),
            data_re_in(7) => data_re_in(502),
            data_re_in(8) => data_re_in(566),
            data_re_in(9) => data_re_in(630),
            data_re_in(10) => data_re_in(694),
            data_re_in(11) => data_re_in(758),
            data_re_in(12) => data_re_in(822),
            data_re_in(13) => data_re_in(886),
            data_re_in(14) => data_re_in(950),
            data_re_in(15) => data_re_in(1014),
            data_re_in(16) => data_re_in(1078),
            data_re_in(17) => data_re_in(1142),
            data_re_in(18) => data_re_in(1206),
            data_re_in(19) => data_re_in(1270),
            data_re_in(20) => data_re_in(1334),
            data_re_in(21) => data_re_in(1398),
            data_re_in(22) => data_re_in(1462),
            data_re_in(23) => data_re_in(1526),
            data_re_in(24) => data_re_in(1590),
            data_re_in(25) => data_re_in(1654),
            data_re_in(26) => data_re_in(1718),
            data_re_in(27) => data_re_in(1782),
            data_re_in(28) => data_re_in(1846),
            data_re_in(29) => data_re_in(1910),
            data_re_in(30) => data_re_in(1974),
            data_re_in(31) => data_re_in(2038),
            data_im_in(0) => data_im_in(54),
            data_im_in(1) => data_im_in(118),
            data_im_in(2) => data_im_in(182),
            data_im_in(3) => data_im_in(246),
            data_im_in(4) => data_im_in(310),
            data_im_in(5) => data_im_in(374),
            data_im_in(6) => data_im_in(438),
            data_im_in(7) => data_im_in(502),
            data_im_in(8) => data_im_in(566),
            data_im_in(9) => data_im_in(630),
            data_im_in(10) => data_im_in(694),
            data_im_in(11) => data_im_in(758),
            data_im_in(12) => data_im_in(822),
            data_im_in(13) => data_im_in(886),
            data_im_in(14) => data_im_in(950),
            data_im_in(15) => data_im_in(1014),
            data_im_in(16) => data_im_in(1078),
            data_im_in(17) => data_im_in(1142),
            data_im_in(18) => data_im_in(1206),
            data_im_in(19) => data_im_in(1270),
            data_im_in(20) => data_im_in(1334),
            data_im_in(21) => data_im_in(1398),
            data_im_in(22) => data_im_in(1462),
            data_im_in(23) => data_im_in(1526),
            data_im_in(24) => data_im_in(1590),
            data_im_in(25) => data_im_in(1654),
            data_im_in(26) => data_im_in(1718),
            data_im_in(27) => data_im_in(1782),
            data_im_in(28) => data_im_in(1846),
            data_im_in(29) => data_im_in(1910),
            data_im_in(30) => data_im_in(1974),
            data_im_in(31) => data_im_in(2038),
            data_re_out(0) => first_stage_re_out(54),
            data_re_out(1) => first_stage_re_out(118),
            data_re_out(2) => first_stage_re_out(182),
            data_re_out(3) => first_stage_re_out(246),
            data_re_out(4) => first_stage_re_out(310),
            data_re_out(5) => first_stage_re_out(374),
            data_re_out(6) => first_stage_re_out(438),
            data_re_out(7) => first_stage_re_out(502),
            data_re_out(8) => first_stage_re_out(566),
            data_re_out(9) => first_stage_re_out(630),
            data_re_out(10) => first_stage_re_out(694),
            data_re_out(11) => first_stage_re_out(758),
            data_re_out(12) => first_stage_re_out(822),
            data_re_out(13) => first_stage_re_out(886),
            data_re_out(14) => first_stage_re_out(950),
            data_re_out(15) => first_stage_re_out(1014),
            data_re_out(16) => first_stage_re_out(1078),
            data_re_out(17) => first_stage_re_out(1142),
            data_re_out(18) => first_stage_re_out(1206),
            data_re_out(19) => first_stage_re_out(1270),
            data_re_out(20) => first_stage_re_out(1334),
            data_re_out(21) => first_stage_re_out(1398),
            data_re_out(22) => first_stage_re_out(1462),
            data_re_out(23) => first_stage_re_out(1526),
            data_re_out(24) => first_stage_re_out(1590),
            data_re_out(25) => first_stage_re_out(1654),
            data_re_out(26) => first_stage_re_out(1718),
            data_re_out(27) => first_stage_re_out(1782),
            data_re_out(28) => first_stage_re_out(1846),
            data_re_out(29) => first_stage_re_out(1910),
            data_re_out(30) => first_stage_re_out(1974),
            data_re_out(31) => first_stage_re_out(2038),
            data_im_out(0) => first_stage_im_out(54),
            data_im_out(1) => first_stage_im_out(118),
            data_im_out(2) => first_stage_im_out(182),
            data_im_out(3) => first_stage_im_out(246),
            data_im_out(4) => first_stage_im_out(310),
            data_im_out(5) => first_stage_im_out(374),
            data_im_out(6) => first_stage_im_out(438),
            data_im_out(7) => first_stage_im_out(502),
            data_im_out(8) => first_stage_im_out(566),
            data_im_out(9) => first_stage_im_out(630),
            data_im_out(10) => first_stage_im_out(694),
            data_im_out(11) => first_stage_im_out(758),
            data_im_out(12) => first_stage_im_out(822),
            data_im_out(13) => first_stage_im_out(886),
            data_im_out(14) => first_stage_im_out(950),
            data_im_out(15) => first_stage_im_out(1014),
            data_im_out(16) => first_stage_im_out(1078),
            data_im_out(17) => first_stage_im_out(1142),
            data_im_out(18) => first_stage_im_out(1206),
            data_im_out(19) => first_stage_im_out(1270),
            data_im_out(20) => first_stage_im_out(1334),
            data_im_out(21) => first_stage_im_out(1398),
            data_im_out(22) => first_stage_im_out(1462),
            data_im_out(23) => first_stage_im_out(1526),
            data_im_out(24) => first_stage_im_out(1590),
            data_im_out(25) => first_stage_im_out(1654),
            data_im_out(26) => first_stage_im_out(1718),
            data_im_out(27) => first_stage_im_out(1782),
            data_im_out(28) => first_stage_im_out(1846),
            data_im_out(29) => first_stage_im_out(1910),
            data_im_out(30) => first_stage_im_out(1974),
            data_im_out(31) => first_stage_im_out(2038)
        );

    ULFFT_PT32_55 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(55),
            data_re_in(1) => data_re_in(119),
            data_re_in(2) => data_re_in(183),
            data_re_in(3) => data_re_in(247),
            data_re_in(4) => data_re_in(311),
            data_re_in(5) => data_re_in(375),
            data_re_in(6) => data_re_in(439),
            data_re_in(7) => data_re_in(503),
            data_re_in(8) => data_re_in(567),
            data_re_in(9) => data_re_in(631),
            data_re_in(10) => data_re_in(695),
            data_re_in(11) => data_re_in(759),
            data_re_in(12) => data_re_in(823),
            data_re_in(13) => data_re_in(887),
            data_re_in(14) => data_re_in(951),
            data_re_in(15) => data_re_in(1015),
            data_re_in(16) => data_re_in(1079),
            data_re_in(17) => data_re_in(1143),
            data_re_in(18) => data_re_in(1207),
            data_re_in(19) => data_re_in(1271),
            data_re_in(20) => data_re_in(1335),
            data_re_in(21) => data_re_in(1399),
            data_re_in(22) => data_re_in(1463),
            data_re_in(23) => data_re_in(1527),
            data_re_in(24) => data_re_in(1591),
            data_re_in(25) => data_re_in(1655),
            data_re_in(26) => data_re_in(1719),
            data_re_in(27) => data_re_in(1783),
            data_re_in(28) => data_re_in(1847),
            data_re_in(29) => data_re_in(1911),
            data_re_in(30) => data_re_in(1975),
            data_re_in(31) => data_re_in(2039),
            data_im_in(0) => data_im_in(55),
            data_im_in(1) => data_im_in(119),
            data_im_in(2) => data_im_in(183),
            data_im_in(3) => data_im_in(247),
            data_im_in(4) => data_im_in(311),
            data_im_in(5) => data_im_in(375),
            data_im_in(6) => data_im_in(439),
            data_im_in(7) => data_im_in(503),
            data_im_in(8) => data_im_in(567),
            data_im_in(9) => data_im_in(631),
            data_im_in(10) => data_im_in(695),
            data_im_in(11) => data_im_in(759),
            data_im_in(12) => data_im_in(823),
            data_im_in(13) => data_im_in(887),
            data_im_in(14) => data_im_in(951),
            data_im_in(15) => data_im_in(1015),
            data_im_in(16) => data_im_in(1079),
            data_im_in(17) => data_im_in(1143),
            data_im_in(18) => data_im_in(1207),
            data_im_in(19) => data_im_in(1271),
            data_im_in(20) => data_im_in(1335),
            data_im_in(21) => data_im_in(1399),
            data_im_in(22) => data_im_in(1463),
            data_im_in(23) => data_im_in(1527),
            data_im_in(24) => data_im_in(1591),
            data_im_in(25) => data_im_in(1655),
            data_im_in(26) => data_im_in(1719),
            data_im_in(27) => data_im_in(1783),
            data_im_in(28) => data_im_in(1847),
            data_im_in(29) => data_im_in(1911),
            data_im_in(30) => data_im_in(1975),
            data_im_in(31) => data_im_in(2039),
            data_re_out(0) => first_stage_re_out(55),
            data_re_out(1) => first_stage_re_out(119),
            data_re_out(2) => first_stage_re_out(183),
            data_re_out(3) => first_stage_re_out(247),
            data_re_out(4) => first_stage_re_out(311),
            data_re_out(5) => first_stage_re_out(375),
            data_re_out(6) => first_stage_re_out(439),
            data_re_out(7) => first_stage_re_out(503),
            data_re_out(8) => first_stage_re_out(567),
            data_re_out(9) => first_stage_re_out(631),
            data_re_out(10) => first_stage_re_out(695),
            data_re_out(11) => first_stage_re_out(759),
            data_re_out(12) => first_stage_re_out(823),
            data_re_out(13) => first_stage_re_out(887),
            data_re_out(14) => first_stage_re_out(951),
            data_re_out(15) => first_stage_re_out(1015),
            data_re_out(16) => first_stage_re_out(1079),
            data_re_out(17) => first_stage_re_out(1143),
            data_re_out(18) => first_stage_re_out(1207),
            data_re_out(19) => first_stage_re_out(1271),
            data_re_out(20) => first_stage_re_out(1335),
            data_re_out(21) => first_stage_re_out(1399),
            data_re_out(22) => first_stage_re_out(1463),
            data_re_out(23) => first_stage_re_out(1527),
            data_re_out(24) => first_stage_re_out(1591),
            data_re_out(25) => first_stage_re_out(1655),
            data_re_out(26) => first_stage_re_out(1719),
            data_re_out(27) => first_stage_re_out(1783),
            data_re_out(28) => first_stage_re_out(1847),
            data_re_out(29) => first_stage_re_out(1911),
            data_re_out(30) => first_stage_re_out(1975),
            data_re_out(31) => first_stage_re_out(2039),
            data_im_out(0) => first_stage_im_out(55),
            data_im_out(1) => first_stage_im_out(119),
            data_im_out(2) => first_stage_im_out(183),
            data_im_out(3) => first_stage_im_out(247),
            data_im_out(4) => first_stage_im_out(311),
            data_im_out(5) => first_stage_im_out(375),
            data_im_out(6) => first_stage_im_out(439),
            data_im_out(7) => first_stage_im_out(503),
            data_im_out(8) => first_stage_im_out(567),
            data_im_out(9) => first_stage_im_out(631),
            data_im_out(10) => first_stage_im_out(695),
            data_im_out(11) => first_stage_im_out(759),
            data_im_out(12) => first_stage_im_out(823),
            data_im_out(13) => first_stage_im_out(887),
            data_im_out(14) => first_stage_im_out(951),
            data_im_out(15) => first_stage_im_out(1015),
            data_im_out(16) => first_stage_im_out(1079),
            data_im_out(17) => first_stage_im_out(1143),
            data_im_out(18) => first_stage_im_out(1207),
            data_im_out(19) => first_stage_im_out(1271),
            data_im_out(20) => first_stage_im_out(1335),
            data_im_out(21) => first_stage_im_out(1399),
            data_im_out(22) => first_stage_im_out(1463),
            data_im_out(23) => first_stage_im_out(1527),
            data_im_out(24) => first_stage_im_out(1591),
            data_im_out(25) => first_stage_im_out(1655),
            data_im_out(26) => first_stage_im_out(1719),
            data_im_out(27) => first_stage_im_out(1783),
            data_im_out(28) => first_stage_im_out(1847),
            data_im_out(29) => first_stage_im_out(1911),
            data_im_out(30) => first_stage_im_out(1975),
            data_im_out(31) => first_stage_im_out(2039)
        );

    ULFFT_PT32_56 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(56),
            data_re_in(1) => data_re_in(120),
            data_re_in(2) => data_re_in(184),
            data_re_in(3) => data_re_in(248),
            data_re_in(4) => data_re_in(312),
            data_re_in(5) => data_re_in(376),
            data_re_in(6) => data_re_in(440),
            data_re_in(7) => data_re_in(504),
            data_re_in(8) => data_re_in(568),
            data_re_in(9) => data_re_in(632),
            data_re_in(10) => data_re_in(696),
            data_re_in(11) => data_re_in(760),
            data_re_in(12) => data_re_in(824),
            data_re_in(13) => data_re_in(888),
            data_re_in(14) => data_re_in(952),
            data_re_in(15) => data_re_in(1016),
            data_re_in(16) => data_re_in(1080),
            data_re_in(17) => data_re_in(1144),
            data_re_in(18) => data_re_in(1208),
            data_re_in(19) => data_re_in(1272),
            data_re_in(20) => data_re_in(1336),
            data_re_in(21) => data_re_in(1400),
            data_re_in(22) => data_re_in(1464),
            data_re_in(23) => data_re_in(1528),
            data_re_in(24) => data_re_in(1592),
            data_re_in(25) => data_re_in(1656),
            data_re_in(26) => data_re_in(1720),
            data_re_in(27) => data_re_in(1784),
            data_re_in(28) => data_re_in(1848),
            data_re_in(29) => data_re_in(1912),
            data_re_in(30) => data_re_in(1976),
            data_re_in(31) => data_re_in(2040),
            data_im_in(0) => data_im_in(56),
            data_im_in(1) => data_im_in(120),
            data_im_in(2) => data_im_in(184),
            data_im_in(3) => data_im_in(248),
            data_im_in(4) => data_im_in(312),
            data_im_in(5) => data_im_in(376),
            data_im_in(6) => data_im_in(440),
            data_im_in(7) => data_im_in(504),
            data_im_in(8) => data_im_in(568),
            data_im_in(9) => data_im_in(632),
            data_im_in(10) => data_im_in(696),
            data_im_in(11) => data_im_in(760),
            data_im_in(12) => data_im_in(824),
            data_im_in(13) => data_im_in(888),
            data_im_in(14) => data_im_in(952),
            data_im_in(15) => data_im_in(1016),
            data_im_in(16) => data_im_in(1080),
            data_im_in(17) => data_im_in(1144),
            data_im_in(18) => data_im_in(1208),
            data_im_in(19) => data_im_in(1272),
            data_im_in(20) => data_im_in(1336),
            data_im_in(21) => data_im_in(1400),
            data_im_in(22) => data_im_in(1464),
            data_im_in(23) => data_im_in(1528),
            data_im_in(24) => data_im_in(1592),
            data_im_in(25) => data_im_in(1656),
            data_im_in(26) => data_im_in(1720),
            data_im_in(27) => data_im_in(1784),
            data_im_in(28) => data_im_in(1848),
            data_im_in(29) => data_im_in(1912),
            data_im_in(30) => data_im_in(1976),
            data_im_in(31) => data_im_in(2040),
            data_re_out(0) => first_stage_re_out(56),
            data_re_out(1) => first_stage_re_out(120),
            data_re_out(2) => first_stage_re_out(184),
            data_re_out(3) => first_stage_re_out(248),
            data_re_out(4) => first_stage_re_out(312),
            data_re_out(5) => first_stage_re_out(376),
            data_re_out(6) => first_stage_re_out(440),
            data_re_out(7) => first_stage_re_out(504),
            data_re_out(8) => first_stage_re_out(568),
            data_re_out(9) => first_stage_re_out(632),
            data_re_out(10) => first_stage_re_out(696),
            data_re_out(11) => first_stage_re_out(760),
            data_re_out(12) => first_stage_re_out(824),
            data_re_out(13) => first_stage_re_out(888),
            data_re_out(14) => first_stage_re_out(952),
            data_re_out(15) => first_stage_re_out(1016),
            data_re_out(16) => first_stage_re_out(1080),
            data_re_out(17) => first_stage_re_out(1144),
            data_re_out(18) => first_stage_re_out(1208),
            data_re_out(19) => first_stage_re_out(1272),
            data_re_out(20) => first_stage_re_out(1336),
            data_re_out(21) => first_stage_re_out(1400),
            data_re_out(22) => first_stage_re_out(1464),
            data_re_out(23) => first_stage_re_out(1528),
            data_re_out(24) => first_stage_re_out(1592),
            data_re_out(25) => first_stage_re_out(1656),
            data_re_out(26) => first_stage_re_out(1720),
            data_re_out(27) => first_stage_re_out(1784),
            data_re_out(28) => first_stage_re_out(1848),
            data_re_out(29) => first_stage_re_out(1912),
            data_re_out(30) => first_stage_re_out(1976),
            data_re_out(31) => first_stage_re_out(2040),
            data_im_out(0) => first_stage_im_out(56),
            data_im_out(1) => first_stage_im_out(120),
            data_im_out(2) => first_stage_im_out(184),
            data_im_out(3) => first_stage_im_out(248),
            data_im_out(4) => first_stage_im_out(312),
            data_im_out(5) => first_stage_im_out(376),
            data_im_out(6) => first_stage_im_out(440),
            data_im_out(7) => first_stage_im_out(504),
            data_im_out(8) => first_stage_im_out(568),
            data_im_out(9) => first_stage_im_out(632),
            data_im_out(10) => first_stage_im_out(696),
            data_im_out(11) => first_stage_im_out(760),
            data_im_out(12) => first_stage_im_out(824),
            data_im_out(13) => first_stage_im_out(888),
            data_im_out(14) => first_stage_im_out(952),
            data_im_out(15) => first_stage_im_out(1016),
            data_im_out(16) => first_stage_im_out(1080),
            data_im_out(17) => first_stage_im_out(1144),
            data_im_out(18) => first_stage_im_out(1208),
            data_im_out(19) => first_stage_im_out(1272),
            data_im_out(20) => first_stage_im_out(1336),
            data_im_out(21) => first_stage_im_out(1400),
            data_im_out(22) => first_stage_im_out(1464),
            data_im_out(23) => first_stage_im_out(1528),
            data_im_out(24) => first_stage_im_out(1592),
            data_im_out(25) => first_stage_im_out(1656),
            data_im_out(26) => first_stage_im_out(1720),
            data_im_out(27) => first_stage_im_out(1784),
            data_im_out(28) => first_stage_im_out(1848),
            data_im_out(29) => first_stage_im_out(1912),
            data_im_out(30) => first_stage_im_out(1976),
            data_im_out(31) => first_stage_im_out(2040)
        );

    ULFFT_PT32_57 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(57),
            data_re_in(1) => data_re_in(121),
            data_re_in(2) => data_re_in(185),
            data_re_in(3) => data_re_in(249),
            data_re_in(4) => data_re_in(313),
            data_re_in(5) => data_re_in(377),
            data_re_in(6) => data_re_in(441),
            data_re_in(7) => data_re_in(505),
            data_re_in(8) => data_re_in(569),
            data_re_in(9) => data_re_in(633),
            data_re_in(10) => data_re_in(697),
            data_re_in(11) => data_re_in(761),
            data_re_in(12) => data_re_in(825),
            data_re_in(13) => data_re_in(889),
            data_re_in(14) => data_re_in(953),
            data_re_in(15) => data_re_in(1017),
            data_re_in(16) => data_re_in(1081),
            data_re_in(17) => data_re_in(1145),
            data_re_in(18) => data_re_in(1209),
            data_re_in(19) => data_re_in(1273),
            data_re_in(20) => data_re_in(1337),
            data_re_in(21) => data_re_in(1401),
            data_re_in(22) => data_re_in(1465),
            data_re_in(23) => data_re_in(1529),
            data_re_in(24) => data_re_in(1593),
            data_re_in(25) => data_re_in(1657),
            data_re_in(26) => data_re_in(1721),
            data_re_in(27) => data_re_in(1785),
            data_re_in(28) => data_re_in(1849),
            data_re_in(29) => data_re_in(1913),
            data_re_in(30) => data_re_in(1977),
            data_re_in(31) => data_re_in(2041),
            data_im_in(0) => data_im_in(57),
            data_im_in(1) => data_im_in(121),
            data_im_in(2) => data_im_in(185),
            data_im_in(3) => data_im_in(249),
            data_im_in(4) => data_im_in(313),
            data_im_in(5) => data_im_in(377),
            data_im_in(6) => data_im_in(441),
            data_im_in(7) => data_im_in(505),
            data_im_in(8) => data_im_in(569),
            data_im_in(9) => data_im_in(633),
            data_im_in(10) => data_im_in(697),
            data_im_in(11) => data_im_in(761),
            data_im_in(12) => data_im_in(825),
            data_im_in(13) => data_im_in(889),
            data_im_in(14) => data_im_in(953),
            data_im_in(15) => data_im_in(1017),
            data_im_in(16) => data_im_in(1081),
            data_im_in(17) => data_im_in(1145),
            data_im_in(18) => data_im_in(1209),
            data_im_in(19) => data_im_in(1273),
            data_im_in(20) => data_im_in(1337),
            data_im_in(21) => data_im_in(1401),
            data_im_in(22) => data_im_in(1465),
            data_im_in(23) => data_im_in(1529),
            data_im_in(24) => data_im_in(1593),
            data_im_in(25) => data_im_in(1657),
            data_im_in(26) => data_im_in(1721),
            data_im_in(27) => data_im_in(1785),
            data_im_in(28) => data_im_in(1849),
            data_im_in(29) => data_im_in(1913),
            data_im_in(30) => data_im_in(1977),
            data_im_in(31) => data_im_in(2041),
            data_re_out(0) => first_stage_re_out(57),
            data_re_out(1) => first_stage_re_out(121),
            data_re_out(2) => first_stage_re_out(185),
            data_re_out(3) => first_stage_re_out(249),
            data_re_out(4) => first_stage_re_out(313),
            data_re_out(5) => first_stage_re_out(377),
            data_re_out(6) => first_stage_re_out(441),
            data_re_out(7) => first_stage_re_out(505),
            data_re_out(8) => first_stage_re_out(569),
            data_re_out(9) => first_stage_re_out(633),
            data_re_out(10) => first_stage_re_out(697),
            data_re_out(11) => first_stage_re_out(761),
            data_re_out(12) => first_stage_re_out(825),
            data_re_out(13) => first_stage_re_out(889),
            data_re_out(14) => first_stage_re_out(953),
            data_re_out(15) => first_stage_re_out(1017),
            data_re_out(16) => first_stage_re_out(1081),
            data_re_out(17) => first_stage_re_out(1145),
            data_re_out(18) => first_stage_re_out(1209),
            data_re_out(19) => first_stage_re_out(1273),
            data_re_out(20) => first_stage_re_out(1337),
            data_re_out(21) => first_stage_re_out(1401),
            data_re_out(22) => first_stage_re_out(1465),
            data_re_out(23) => first_stage_re_out(1529),
            data_re_out(24) => first_stage_re_out(1593),
            data_re_out(25) => first_stage_re_out(1657),
            data_re_out(26) => first_stage_re_out(1721),
            data_re_out(27) => first_stage_re_out(1785),
            data_re_out(28) => first_stage_re_out(1849),
            data_re_out(29) => first_stage_re_out(1913),
            data_re_out(30) => first_stage_re_out(1977),
            data_re_out(31) => first_stage_re_out(2041),
            data_im_out(0) => first_stage_im_out(57),
            data_im_out(1) => first_stage_im_out(121),
            data_im_out(2) => first_stage_im_out(185),
            data_im_out(3) => first_stage_im_out(249),
            data_im_out(4) => first_stage_im_out(313),
            data_im_out(5) => first_stage_im_out(377),
            data_im_out(6) => first_stage_im_out(441),
            data_im_out(7) => first_stage_im_out(505),
            data_im_out(8) => first_stage_im_out(569),
            data_im_out(9) => first_stage_im_out(633),
            data_im_out(10) => first_stage_im_out(697),
            data_im_out(11) => first_stage_im_out(761),
            data_im_out(12) => first_stage_im_out(825),
            data_im_out(13) => first_stage_im_out(889),
            data_im_out(14) => first_stage_im_out(953),
            data_im_out(15) => first_stage_im_out(1017),
            data_im_out(16) => first_stage_im_out(1081),
            data_im_out(17) => first_stage_im_out(1145),
            data_im_out(18) => first_stage_im_out(1209),
            data_im_out(19) => first_stage_im_out(1273),
            data_im_out(20) => first_stage_im_out(1337),
            data_im_out(21) => first_stage_im_out(1401),
            data_im_out(22) => first_stage_im_out(1465),
            data_im_out(23) => first_stage_im_out(1529),
            data_im_out(24) => first_stage_im_out(1593),
            data_im_out(25) => first_stage_im_out(1657),
            data_im_out(26) => first_stage_im_out(1721),
            data_im_out(27) => first_stage_im_out(1785),
            data_im_out(28) => first_stage_im_out(1849),
            data_im_out(29) => first_stage_im_out(1913),
            data_im_out(30) => first_stage_im_out(1977),
            data_im_out(31) => first_stage_im_out(2041)
        );

    ULFFT_PT32_58 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(58),
            data_re_in(1) => data_re_in(122),
            data_re_in(2) => data_re_in(186),
            data_re_in(3) => data_re_in(250),
            data_re_in(4) => data_re_in(314),
            data_re_in(5) => data_re_in(378),
            data_re_in(6) => data_re_in(442),
            data_re_in(7) => data_re_in(506),
            data_re_in(8) => data_re_in(570),
            data_re_in(9) => data_re_in(634),
            data_re_in(10) => data_re_in(698),
            data_re_in(11) => data_re_in(762),
            data_re_in(12) => data_re_in(826),
            data_re_in(13) => data_re_in(890),
            data_re_in(14) => data_re_in(954),
            data_re_in(15) => data_re_in(1018),
            data_re_in(16) => data_re_in(1082),
            data_re_in(17) => data_re_in(1146),
            data_re_in(18) => data_re_in(1210),
            data_re_in(19) => data_re_in(1274),
            data_re_in(20) => data_re_in(1338),
            data_re_in(21) => data_re_in(1402),
            data_re_in(22) => data_re_in(1466),
            data_re_in(23) => data_re_in(1530),
            data_re_in(24) => data_re_in(1594),
            data_re_in(25) => data_re_in(1658),
            data_re_in(26) => data_re_in(1722),
            data_re_in(27) => data_re_in(1786),
            data_re_in(28) => data_re_in(1850),
            data_re_in(29) => data_re_in(1914),
            data_re_in(30) => data_re_in(1978),
            data_re_in(31) => data_re_in(2042),
            data_im_in(0) => data_im_in(58),
            data_im_in(1) => data_im_in(122),
            data_im_in(2) => data_im_in(186),
            data_im_in(3) => data_im_in(250),
            data_im_in(4) => data_im_in(314),
            data_im_in(5) => data_im_in(378),
            data_im_in(6) => data_im_in(442),
            data_im_in(7) => data_im_in(506),
            data_im_in(8) => data_im_in(570),
            data_im_in(9) => data_im_in(634),
            data_im_in(10) => data_im_in(698),
            data_im_in(11) => data_im_in(762),
            data_im_in(12) => data_im_in(826),
            data_im_in(13) => data_im_in(890),
            data_im_in(14) => data_im_in(954),
            data_im_in(15) => data_im_in(1018),
            data_im_in(16) => data_im_in(1082),
            data_im_in(17) => data_im_in(1146),
            data_im_in(18) => data_im_in(1210),
            data_im_in(19) => data_im_in(1274),
            data_im_in(20) => data_im_in(1338),
            data_im_in(21) => data_im_in(1402),
            data_im_in(22) => data_im_in(1466),
            data_im_in(23) => data_im_in(1530),
            data_im_in(24) => data_im_in(1594),
            data_im_in(25) => data_im_in(1658),
            data_im_in(26) => data_im_in(1722),
            data_im_in(27) => data_im_in(1786),
            data_im_in(28) => data_im_in(1850),
            data_im_in(29) => data_im_in(1914),
            data_im_in(30) => data_im_in(1978),
            data_im_in(31) => data_im_in(2042),
            data_re_out(0) => first_stage_re_out(58),
            data_re_out(1) => first_stage_re_out(122),
            data_re_out(2) => first_stage_re_out(186),
            data_re_out(3) => first_stage_re_out(250),
            data_re_out(4) => first_stage_re_out(314),
            data_re_out(5) => first_stage_re_out(378),
            data_re_out(6) => first_stage_re_out(442),
            data_re_out(7) => first_stage_re_out(506),
            data_re_out(8) => first_stage_re_out(570),
            data_re_out(9) => first_stage_re_out(634),
            data_re_out(10) => first_stage_re_out(698),
            data_re_out(11) => first_stage_re_out(762),
            data_re_out(12) => first_stage_re_out(826),
            data_re_out(13) => first_stage_re_out(890),
            data_re_out(14) => first_stage_re_out(954),
            data_re_out(15) => first_stage_re_out(1018),
            data_re_out(16) => first_stage_re_out(1082),
            data_re_out(17) => first_stage_re_out(1146),
            data_re_out(18) => first_stage_re_out(1210),
            data_re_out(19) => first_stage_re_out(1274),
            data_re_out(20) => first_stage_re_out(1338),
            data_re_out(21) => first_stage_re_out(1402),
            data_re_out(22) => first_stage_re_out(1466),
            data_re_out(23) => first_stage_re_out(1530),
            data_re_out(24) => first_stage_re_out(1594),
            data_re_out(25) => first_stage_re_out(1658),
            data_re_out(26) => first_stage_re_out(1722),
            data_re_out(27) => first_stage_re_out(1786),
            data_re_out(28) => first_stage_re_out(1850),
            data_re_out(29) => first_stage_re_out(1914),
            data_re_out(30) => first_stage_re_out(1978),
            data_re_out(31) => first_stage_re_out(2042),
            data_im_out(0) => first_stage_im_out(58),
            data_im_out(1) => first_stage_im_out(122),
            data_im_out(2) => first_stage_im_out(186),
            data_im_out(3) => first_stage_im_out(250),
            data_im_out(4) => first_stage_im_out(314),
            data_im_out(5) => first_stage_im_out(378),
            data_im_out(6) => first_stage_im_out(442),
            data_im_out(7) => first_stage_im_out(506),
            data_im_out(8) => first_stage_im_out(570),
            data_im_out(9) => first_stage_im_out(634),
            data_im_out(10) => first_stage_im_out(698),
            data_im_out(11) => first_stage_im_out(762),
            data_im_out(12) => first_stage_im_out(826),
            data_im_out(13) => first_stage_im_out(890),
            data_im_out(14) => first_stage_im_out(954),
            data_im_out(15) => first_stage_im_out(1018),
            data_im_out(16) => first_stage_im_out(1082),
            data_im_out(17) => first_stage_im_out(1146),
            data_im_out(18) => first_stage_im_out(1210),
            data_im_out(19) => first_stage_im_out(1274),
            data_im_out(20) => first_stage_im_out(1338),
            data_im_out(21) => first_stage_im_out(1402),
            data_im_out(22) => first_stage_im_out(1466),
            data_im_out(23) => first_stage_im_out(1530),
            data_im_out(24) => first_stage_im_out(1594),
            data_im_out(25) => first_stage_im_out(1658),
            data_im_out(26) => first_stage_im_out(1722),
            data_im_out(27) => first_stage_im_out(1786),
            data_im_out(28) => first_stage_im_out(1850),
            data_im_out(29) => first_stage_im_out(1914),
            data_im_out(30) => first_stage_im_out(1978),
            data_im_out(31) => first_stage_im_out(2042)
        );

    ULFFT_PT32_59 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(59),
            data_re_in(1) => data_re_in(123),
            data_re_in(2) => data_re_in(187),
            data_re_in(3) => data_re_in(251),
            data_re_in(4) => data_re_in(315),
            data_re_in(5) => data_re_in(379),
            data_re_in(6) => data_re_in(443),
            data_re_in(7) => data_re_in(507),
            data_re_in(8) => data_re_in(571),
            data_re_in(9) => data_re_in(635),
            data_re_in(10) => data_re_in(699),
            data_re_in(11) => data_re_in(763),
            data_re_in(12) => data_re_in(827),
            data_re_in(13) => data_re_in(891),
            data_re_in(14) => data_re_in(955),
            data_re_in(15) => data_re_in(1019),
            data_re_in(16) => data_re_in(1083),
            data_re_in(17) => data_re_in(1147),
            data_re_in(18) => data_re_in(1211),
            data_re_in(19) => data_re_in(1275),
            data_re_in(20) => data_re_in(1339),
            data_re_in(21) => data_re_in(1403),
            data_re_in(22) => data_re_in(1467),
            data_re_in(23) => data_re_in(1531),
            data_re_in(24) => data_re_in(1595),
            data_re_in(25) => data_re_in(1659),
            data_re_in(26) => data_re_in(1723),
            data_re_in(27) => data_re_in(1787),
            data_re_in(28) => data_re_in(1851),
            data_re_in(29) => data_re_in(1915),
            data_re_in(30) => data_re_in(1979),
            data_re_in(31) => data_re_in(2043),
            data_im_in(0) => data_im_in(59),
            data_im_in(1) => data_im_in(123),
            data_im_in(2) => data_im_in(187),
            data_im_in(3) => data_im_in(251),
            data_im_in(4) => data_im_in(315),
            data_im_in(5) => data_im_in(379),
            data_im_in(6) => data_im_in(443),
            data_im_in(7) => data_im_in(507),
            data_im_in(8) => data_im_in(571),
            data_im_in(9) => data_im_in(635),
            data_im_in(10) => data_im_in(699),
            data_im_in(11) => data_im_in(763),
            data_im_in(12) => data_im_in(827),
            data_im_in(13) => data_im_in(891),
            data_im_in(14) => data_im_in(955),
            data_im_in(15) => data_im_in(1019),
            data_im_in(16) => data_im_in(1083),
            data_im_in(17) => data_im_in(1147),
            data_im_in(18) => data_im_in(1211),
            data_im_in(19) => data_im_in(1275),
            data_im_in(20) => data_im_in(1339),
            data_im_in(21) => data_im_in(1403),
            data_im_in(22) => data_im_in(1467),
            data_im_in(23) => data_im_in(1531),
            data_im_in(24) => data_im_in(1595),
            data_im_in(25) => data_im_in(1659),
            data_im_in(26) => data_im_in(1723),
            data_im_in(27) => data_im_in(1787),
            data_im_in(28) => data_im_in(1851),
            data_im_in(29) => data_im_in(1915),
            data_im_in(30) => data_im_in(1979),
            data_im_in(31) => data_im_in(2043),
            data_re_out(0) => first_stage_re_out(59),
            data_re_out(1) => first_stage_re_out(123),
            data_re_out(2) => first_stage_re_out(187),
            data_re_out(3) => first_stage_re_out(251),
            data_re_out(4) => first_stage_re_out(315),
            data_re_out(5) => first_stage_re_out(379),
            data_re_out(6) => first_stage_re_out(443),
            data_re_out(7) => first_stage_re_out(507),
            data_re_out(8) => first_stage_re_out(571),
            data_re_out(9) => first_stage_re_out(635),
            data_re_out(10) => first_stage_re_out(699),
            data_re_out(11) => first_stage_re_out(763),
            data_re_out(12) => first_stage_re_out(827),
            data_re_out(13) => first_stage_re_out(891),
            data_re_out(14) => first_stage_re_out(955),
            data_re_out(15) => first_stage_re_out(1019),
            data_re_out(16) => first_stage_re_out(1083),
            data_re_out(17) => first_stage_re_out(1147),
            data_re_out(18) => first_stage_re_out(1211),
            data_re_out(19) => first_stage_re_out(1275),
            data_re_out(20) => first_stage_re_out(1339),
            data_re_out(21) => first_stage_re_out(1403),
            data_re_out(22) => first_stage_re_out(1467),
            data_re_out(23) => first_stage_re_out(1531),
            data_re_out(24) => first_stage_re_out(1595),
            data_re_out(25) => first_stage_re_out(1659),
            data_re_out(26) => first_stage_re_out(1723),
            data_re_out(27) => first_stage_re_out(1787),
            data_re_out(28) => first_stage_re_out(1851),
            data_re_out(29) => first_stage_re_out(1915),
            data_re_out(30) => first_stage_re_out(1979),
            data_re_out(31) => first_stage_re_out(2043),
            data_im_out(0) => first_stage_im_out(59),
            data_im_out(1) => first_stage_im_out(123),
            data_im_out(2) => first_stage_im_out(187),
            data_im_out(3) => first_stage_im_out(251),
            data_im_out(4) => first_stage_im_out(315),
            data_im_out(5) => first_stage_im_out(379),
            data_im_out(6) => first_stage_im_out(443),
            data_im_out(7) => first_stage_im_out(507),
            data_im_out(8) => first_stage_im_out(571),
            data_im_out(9) => first_stage_im_out(635),
            data_im_out(10) => first_stage_im_out(699),
            data_im_out(11) => first_stage_im_out(763),
            data_im_out(12) => first_stage_im_out(827),
            data_im_out(13) => first_stage_im_out(891),
            data_im_out(14) => first_stage_im_out(955),
            data_im_out(15) => first_stage_im_out(1019),
            data_im_out(16) => first_stage_im_out(1083),
            data_im_out(17) => first_stage_im_out(1147),
            data_im_out(18) => first_stage_im_out(1211),
            data_im_out(19) => first_stage_im_out(1275),
            data_im_out(20) => first_stage_im_out(1339),
            data_im_out(21) => first_stage_im_out(1403),
            data_im_out(22) => first_stage_im_out(1467),
            data_im_out(23) => first_stage_im_out(1531),
            data_im_out(24) => first_stage_im_out(1595),
            data_im_out(25) => first_stage_im_out(1659),
            data_im_out(26) => first_stage_im_out(1723),
            data_im_out(27) => first_stage_im_out(1787),
            data_im_out(28) => first_stage_im_out(1851),
            data_im_out(29) => first_stage_im_out(1915),
            data_im_out(30) => first_stage_im_out(1979),
            data_im_out(31) => first_stage_im_out(2043)
        );

    ULFFT_PT32_60 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(60),
            data_re_in(1) => data_re_in(124),
            data_re_in(2) => data_re_in(188),
            data_re_in(3) => data_re_in(252),
            data_re_in(4) => data_re_in(316),
            data_re_in(5) => data_re_in(380),
            data_re_in(6) => data_re_in(444),
            data_re_in(7) => data_re_in(508),
            data_re_in(8) => data_re_in(572),
            data_re_in(9) => data_re_in(636),
            data_re_in(10) => data_re_in(700),
            data_re_in(11) => data_re_in(764),
            data_re_in(12) => data_re_in(828),
            data_re_in(13) => data_re_in(892),
            data_re_in(14) => data_re_in(956),
            data_re_in(15) => data_re_in(1020),
            data_re_in(16) => data_re_in(1084),
            data_re_in(17) => data_re_in(1148),
            data_re_in(18) => data_re_in(1212),
            data_re_in(19) => data_re_in(1276),
            data_re_in(20) => data_re_in(1340),
            data_re_in(21) => data_re_in(1404),
            data_re_in(22) => data_re_in(1468),
            data_re_in(23) => data_re_in(1532),
            data_re_in(24) => data_re_in(1596),
            data_re_in(25) => data_re_in(1660),
            data_re_in(26) => data_re_in(1724),
            data_re_in(27) => data_re_in(1788),
            data_re_in(28) => data_re_in(1852),
            data_re_in(29) => data_re_in(1916),
            data_re_in(30) => data_re_in(1980),
            data_re_in(31) => data_re_in(2044),
            data_im_in(0) => data_im_in(60),
            data_im_in(1) => data_im_in(124),
            data_im_in(2) => data_im_in(188),
            data_im_in(3) => data_im_in(252),
            data_im_in(4) => data_im_in(316),
            data_im_in(5) => data_im_in(380),
            data_im_in(6) => data_im_in(444),
            data_im_in(7) => data_im_in(508),
            data_im_in(8) => data_im_in(572),
            data_im_in(9) => data_im_in(636),
            data_im_in(10) => data_im_in(700),
            data_im_in(11) => data_im_in(764),
            data_im_in(12) => data_im_in(828),
            data_im_in(13) => data_im_in(892),
            data_im_in(14) => data_im_in(956),
            data_im_in(15) => data_im_in(1020),
            data_im_in(16) => data_im_in(1084),
            data_im_in(17) => data_im_in(1148),
            data_im_in(18) => data_im_in(1212),
            data_im_in(19) => data_im_in(1276),
            data_im_in(20) => data_im_in(1340),
            data_im_in(21) => data_im_in(1404),
            data_im_in(22) => data_im_in(1468),
            data_im_in(23) => data_im_in(1532),
            data_im_in(24) => data_im_in(1596),
            data_im_in(25) => data_im_in(1660),
            data_im_in(26) => data_im_in(1724),
            data_im_in(27) => data_im_in(1788),
            data_im_in(28) => data_im_in(1852),
            data_im_in(29) => data_im_in(1916),
            data_im_in(30) => data_im_in(1980),
            data_im_in(31) => data_im_in(2044),
            data_re_out(0) => first_stage_re_out(60),
            data_re_out(1) => first_stage_re_out(124),
            data_re_out(2) => first_stage_re_out(188),
            data_re_out(3) => first_stage_re_out(252),
            data_re_out(4) => first_stage_re_out(316),
            data_re_out(5) => first_stage_re_out(380),
            data_re_out(6) => first_stage_re_out(444),
            data_re_out(7) => first_stage_re_out(508),
            data_re_out(8) => first_stage_re_out(572),
            data_re_out(9) => first_stage_re_out(636),
            data_re_out(10) => first_stage_re_out(700),
            data_re_out(11) => first_stage_re_out(764),
            data_re_out(12) => first_stage_re_out(828),
            data_re_out(13) => first_stage_re_out(892),
            data_re_out(14) => first_stage_re_out(956),
            data_re_out(15) => first_stage_re_out(1020),
            data_re_out(16) => first_stage_re_out(1084),
            data_re_out(17) => first_stage_re_out(1148),
            data_re_out(18) => first_stage_re_out(1212),
            data_re_out(19) => first_stage_re_out(1276),
            data_re_out(20) => first_stage_re_out(1340),
            data_re_out(21) => first_stage_re_out(1404),
            data_re_out(22) => first_stage_re_out(1468),
            data_re_out(23) => first_stage_re_out(1532),
            data_re_out(24) => first_stage_re_out(1596),
            data_re_out(25) => first_stage_re_out(1660),
            data_re_out(26) => first_stage_re_out(1724),
            data_re_out(27) => first_stage_re_out(1788),
            data_re_out(28) => first_stage_re_out(1852),
            data_re_out(29) => first_stage_re_out(1916),
            data_re_out(30) => first_stage_re_out(1980),
            data_re_out(31) => first_stage_re_out(2044),
            data_im_out(0) => first_stage_im_out(60),
            data_im_out(1) => first_stage_im_out(124),
            data_im_out(2) => first_stage_im_out(188),
            data_im_out(3) => first_stage_im_out(252),
            data_im_out(4) => first_stage_im_out(316),
            data_im_out(5) => first_stage_im_out(380),
            data_im_out(6) => first_stage_im_out(444),
            data_im_out(7) => first_stage_im_out(508),
            data_im_out(8) => first_stage_im_out(572),
            data_im_out(9) => first_stage_im_out(636),
            data_im_out(10) => first_stage_im_out(700),
            data_im_out(11) => first_stage_im_out(764),
            data_im_out(12) => first_stage_im_out(828),
            data_im_out(13) => first_stage_im_out(892),
            data_im_out(14) => first_stage_im_out(956),
            data_im_out(15) => first_stage_im_out(1020),
            data_im_out(16) => first_stage_im_out(1084),
            data_im_out(17) => first_stage_im_out(1148),
            data_im_out(18) => first_stage_im_out(1212),
            data_im_out(19) => first_stage_im_out(1276),
            data_im_out(20) => first_stage_im_out(1340),
            data_im_out(21) => first_stage_im_out(1404),
            data_im_out(22) => first_stage_im_out(1468),
            data_im_out(23) => first_stage_im_out(1532),
            data_im_out(24) => first_stage_im_out(1596),
            data_im_out(25) => first_stage_im_out(1660),
            data_im_out(26) => first_stage_im_out(1724),
            data_im_out(27) => first_stage_im_out(1788),
            data_im_out(28) => first_stage_im_out(1852),
            data_im_out(29) => first_stage_im_out(1916),
            data_im_out(30) => first_stage_im_out(1980),
            data_im_out(31) => first_stage_im_out(2044)
        );

    ULFFT_PT32_61 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(61),
            data_re_in(1) => data_re_in(125),
            data_re_in(2) => data_re_in(189),
            data_re_in(3) => data_re_in(253),
            data_re_in(4) => data_re_in(317),
            data_re_in(5) => data_re_in(381),
            data_re_in(6) => data_re_in(445),
            data_re_in(7) => data_re_in(509),
            data_re_in(8) => data_re_in(573),
            data_re_in(9) => data_re_in(637),
            data_re_in(10) => data_re_in(701),
            data_re_in(11) => data_re_in(765),
            data_re_in(12) => data_re_in(829),
            data_re_in(13) => data_re_in(893),
            data_re_in(14) => data_re_in(957),
            data_re_in(15) => data_re_in(1021),
            data_re_in(16) => data_re_in(1085),
            data_re_in(17) => data_re_in(1149),
            data_re_in(18) => data_re_in(1213),
            data_re_in(19) => data_re_in(1277),
            data_re_in(20) => data_re_in(1341),
            data_re_in(21) => data_re_in(1405),
            data_re_in(22) => data_re_in(1469),
            data_re_in(23) => data_re_in(1533),
            data_re_in(24) => data_re_in(1597),
            data_re_in(25) => data_re_in(1661),
            data_re_in(26) => data_re_in(1725),
            data_re_in(27) => data_re_in(1789),
            data_re_in(28) => data_re_in(1853),
            data_re_in(29) => data_re_in(1917),
            data_re_in(30) => data_re_in(1981),
            data_re_in(31) => data_re_in(2045),
            data_im_in(0) => data_im_in(61),
            data_im_in(1) => data_im_in(125),
            data_im_in(2) => data_im_in(189),
            data_im_in(3) => data_im_in(253),
            data_im_in(4) => data_im_in(317),
            data_im_in(5) => data_im_in(381),
            data_im_in(6) => data_im_in(445),
            data_im_in(7) => data_im_in(509),
            data_im_in(8) => data_im_in(573),
            data_im_in(9) => data_im_in(637),
            data_im_in(10) => data_im_in(701),
            data_im_in(11) => data_im_in(765),
            data_im_in(12) => data_im_in(829),
            data_im_in(13) => data_im_in(893),
            data_im_in(14) => data_im_in(957),
            data_im_in(15) => data_im_in(1021),
            data_im_in(16) => data_im_in(1085),
            data_im_in(17) => data_im_in(1149),
            data_im_in(18) => data_im_in(1213),
            data_im_in(19) => data_im_in(1277),
            data_im_in(20) => data_im_in(1341),
            data_im_in(21) => data_im_in(1405),
            data_im_in(22) => data_im_in(1469),
            data_im_in(23) => data_im_in(1533),
            data_im_in(24) => data_im_in(1597),
            data_im_in(25) => data_im_in(1661),
            data_im_in(26) => data_im_in(1725),
            data_im_in(27) => data_im_in(1789),
            data_im_in(28) => data_im_in(1853),
            data_im_in(29) => data_im_in(1917),
            data_im_in(30) => data_im_in(1981),
            data_im_in(31) => data_im_in(2045),
            data_re_out(0) => first_stage_re_out(61),
            data_re_out(1) => first_stage_re_out(125),
            data_re_out(2) => first_stage_re_out(189),
            data_re_out(3) => first_stage_re_out(253),
            data_re_out(4) => first_stage_re_out(317),
            data_re_out(5) => first_stage_re_out(381),
            data_re_out(6) => first_stage_re_out(445),
            data_re_out(7) => first_stage_re_out(509),
            data_re_out(8) => first_stage_re_out(573),
            data_re_out(9) => first_stage_re_out(637),
            data_re_out(10) => first_stage_re_out(701),
            data_re_out(11) => first_stage_re_out(765),
            data_re_out(12) => first_stage_re_out(829),
            data_re_out(13) => first_stage_re_out(893),
            data_re_out(14) => first_stage_re_out(957),
            data_re_out(15) => first_stage_re_out(1021),
            data_re_out(16) => first_stage_re_out(1085),
            data_re_out(17) => first_stage_re_out(1149),
            data_re_out(18) => first_stage_re_out(1213),
            data_re_out(19) => first_stage_re_out(1277),
            data_re_out(20) => first_stage_re_out(1341),
            data_re_out(21) => first_stage_re_out(1405),
            data_re_out(22) => first_stage_re_out(1469),
            data_re_out(23) => first_stage_re_out(1533),
            data_re_out(24) => first_stage_re_out(1597),
            data_re_out(25) => first_stage_re_out(1661),
            data_re_out(26) => first_stage_re_out(1725),
            data_re_out(27) => first_stage_re_out(1789),
            data_re_out(28) => first_stage_re_out(1853),
            data_re_out(29) => first_stage_re_out(1917),
            data_re_out(30) => first_stage_re_out(1981),
            data_re_out(31) => first_stage_re_out(2045),
            data_im_out(0) => first_stage_im_out(61),
            data_im_out(1) => first_stage_im_out(125),
            data_im_out(2) => first_stage_im_out(189),
            data_im_out(3) => first_stage_im_out(253),
            data_im_out(4) => first_stage_im_out(317),
            data_im_out(5) => first_stage_im_out(381),
            data_im_out(6) => first_stage_im_out(445),
            data_im_out(7) => first_stage_im_out(509),
            data_im_out(8) => first_stage_im_out(573),
            data_im_out(9) => first_stage_im_out(637),
            data_im_out(10) => first_stage_im_out(701),
            data_im_out(11) => first_stage_im_out(765),
            data_im_out(12) => first_stage_im_out(829),
            data_im_out(13) => first_stage_im_out(893),
            data_im_out(14) => first_stage_im_out(957),
            data_im_out(15) => first_stage_im_out(1021),
            data_im_out(16) => first_stage_im_out(1085),
            data_im_out(17) => first_stage_im_out(1149),
            data_im_out(18) => first_stage_im_out(1213),
            data_im_out(19) => first_stage_im_out(1277),
            data_im_out(20) => first_stage_im_out(1341),
            data_im_out(21) => first_stage_im_out(1405),
            data_im_out(22) => first_stage_im_out(1469),
            data_im_out(23) => first_stage_im_out(1533),
            data_im_out(24) => first_stage_im_out(1597),
            data_im_out(25) => first_stage_im_out(1661),
            data_im_out(26) => first_stage_im_out(1725),
            data_im_out(27) => first_stage_im_out(1789),
            data_im_out(28) => first_stage_im_out(1853),
            data_im_out(29) => first_stage_im_out(1917),
            data_im_out(30) => first_stage_im_out(1981),
            data_im_out(31) => first_stage_im_out(2045)
        );

    ULFFT_PT32_62 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(62),
            data_re_in(1) => data_re_in(126),
            data_re_in(2) => data_re_in(190),
            data_re_in(3) => data_re_in(254),
            data_re_in(4) => data_re_in(318),
            data_re_in(5) => data_re_in(382),
            data_re_in(6) => data_re_in(446),
            data_re_in(7) => data_re_in(510),
            data_re_in(8) => data_re_in(574),
            data_re_in(9) => data_re_in(638),
            data_re_in(10) => data_re_in(702),
            data_re_in(11) => data_re_in(766),
            data_re_in(12) => data_re_in(830),
            data_re_in(13) => data_re_in(894),
            data_re_in(14) => data_re_in(958),
            data_re_in(15) => data_re_in(1022),
            data_re_in(16) => data_re_in(1086),
            data_re_in(17) => data_re_in(1150),
            data_re_in(18) => data_re_in(1214),
            data_re_in(19) => data_re_in(1278),
            data_re_in(20) => data_re_in(1342),
            data_re_in(21) => data_re_in(1406),
            data_re_in(22) => data_re_in(1470),
            data_re_in(23) => data_re_in(1534),
            data_re_in(24) => data_re_in(1598),
            data_re_in(25) => data_re_in(1662),
            data_re_in(26) => data_re_in(1726),
            data_re_in(27) => data_re_in(1790),
            data_re_in(28) => data_re_in(1854),
            data_re_in(29) => data_re_in(1918),
            data_re_in(30) => data_re_in(1982),
            data_re_in(31) => data_re_in(2046),
            data_im_in(0) => data_im_in(62),
            data_im_in(1) => data_im_in(126),
            data_im_in(2) => data_im_in(190),
            data_im_in(3) => data_im_in(254),
            data_im_in(4) => data_im_in(318),
            data_im_in(5) => data_im_in(382),
            data_im_in(6) => data_im_in(446),
            data_im_in(7) => data_im_in(510),
            data_im_in(8) => data_im_in(574),
            data_im_in(9) => data_im_in(638),
            data_im_in(10) => data_im_in(702),
            data_im_in(11) => data_im_in(766),
            data_im_in(12) => data_im_in(830),
            data_im_in(13) => data_im_in(894),
            data_im_in(14) => data_im_in(958),
            data_im_in(15) => data_im_in(1022),
            data_im_in(16) => data_im_in(1086),
            data_im_in(17) => data_im_in(1150),
            data_im_in(18) => data_im_in(1214),
            data_im_in(19) => data_im_in(1278),
            data_im_in(20) => data_im_in(1342),
            data_im_in(21) => data_im_in(1406),
            data_im_in(22) => data_im_in(1470),
            data_im_in(23) => data_im_in(1534),
            data_im_in(24) => data_im_in(1598),
            data_im_in(25) => data_im_in(1662),
            data_im_in(26) => data_im_in(1726),
            data_im_in(27) => data_im_in(1790),
            data_im_in(28) => data_im_in(1854),
            data_im_in(29) => data_im_in(1918),
            data_im_in(30) => data_im_in(1982),
            data_im_in(31) => data_im_in(2046),
            data_re_out(0) => first_stage_re_out(62),
            data_re_out(1) => first_stage_re_out(126),
            data_re_out(2) => first_stage_re_out(190),
            data_re_out(3) => first_stage_re_out(254),
            data_re_out(4) => first_stage_re_out(318),
            data_re_out(5) => first_stage_re_out(382),
            data_re_out(6) => first_stage_re_out(446),
            data_re_out(7) => first_stage_re_out(510),
            data_re_out(8) => first_stage_re_out(574),
            data_re_out(9) => first_stage_re_out(638),
            data_re_out(10) => first_stage_re_out(702),
            data_re_out(11) => first_stage_re_out(766),
            data_re_out(12) => first_stage_re_out(830),
            data_re_out(13) => first_stage_re_out(894),
            data_re_out(14) => first_stage_re_out(958),
            data_re_out(15) => first_stage_re_out(1022),
            data_re_out(16) => first_stage_re_out(1086),
            data_re_out(17) => first_stage_re_out(1150),
            data_re_out(18) => first_stage_re_out(1214),
            data_re_out(19) => first_stage_re_out(1278),
            data_re_out(20) => first_stage_re_out(1342),
            data_re_out(21) => first_stage_re_out(1406),
            data_re_out(22) => first_stage_re_out(1470),
            data_re_out(23) => first_stage_re_out(1534),
            data_re_out(24) => first_stage_re_out(1598),
            data_re_out(25) => first_stage_re_out(1662),
            data_re_out(26) => first_stage_re_out(1726),
            data_re_out(27) => first_stage_re_out(1790),
            data_re_out(28) => first_stage_re_out(1854),
            data_re_out(29) => first_stage_re_out(1918),
            data_re_out(30) => first_stage_re_out(1982),
            data_re_out(31) => first_stage_re_out(2046),
            data_im_out(0) => first_stage_im_out(62),
            data_im_out(1) => first_stage_im_out(126),
            data_im_out(2) => first_stage_im_out(190),
            data_im_out(3) => first_stage_im_out(254),
            data_im_out(4) => first_stage_im_out(318),
            data_im_out(5) => first_stage_im_out(382),
            data_im_out(6) => first_stage_im_out(446),
            data_im_out(7) => first_stage_im_out(510),
            data_im_out(8) => first_stage_im_out(574),
            data_im_out(9) => first_stage_im_out(638),
            data_im_out(10) => first_stage_im_out(702),
            data_im_out(11) => first_stage_im_out(766),
            data_im_out(12) => first_stage_im_out(830),
            data_im_out(13) => first_stage_im_out(894),
            data_im_out(14) => first_stage_im_out(958),
            data_im_out(15) => first_stage_im_out(1022),
            data_im_out(16) => first_stage_im_out(1086),
            data_im_out(17) => first_stage_im_out(1150),
            data_im_out(18) => first_stage_im_out(1214),
            data_im_out(19) => first_stage_im_out(1278),
            data_im_out(20) => first_stage_im_out(1342),
            data_im_out(21) => first_stage_im_out(1406),
            data_im_out(22) => first_stage_im_out(1470),
            data_im_out(23) => first_stage_im_out(1534),
            data_im_out(24) => first_stage_im_out(1598),
            data_im_out(25) => first_stage_im_out(1662),
            data_im_out(26) => first_stage_im_out(1726),
            data_im_out(27) => first_stage_im_out(1790),
            data_im_out(28) => first_stage_im_out(1854),
            data_im_out(29) => first_stage_im_out(1918),
            data_im_out(30) => first_stage_im_out(1982),
            data_im_out(31) => first_stage_im_out(2046)
        );

    ULFFT_PT32_63 : fft_pt32
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass,
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(63),
            data_re_in(1) => data_re_in(127),
            data_re_in(2) => data_re_in(191),
            data_re_in(3) => data_re_in(255),
            data_re_in(4) => data_re_in(319),
            data_re_in(5) => data_re_in(383),
            data_re_in(6) => data_re_in(447),
            data_re_in(7) => data_re_in(511),
            data_re_in(8) => data_re_in(575),
            data_re_in(9) => data_re_in(639),
            data_re_in(10) => data_re_in(703),
            data_re_in(11) => data_re_in(767),
            data_re_in(12) => data_re_in(831),
            data_re_in(13) => data_re_in(895),
            data_re_in(14) => data_re_in(959),
            data_re_in(15) => data_re_in(1023),
            data_re_in(16) => data_re_in(1087),
            data_re_in(17) => data_re_in(1151),
            data_re_in(18) => data_re_in(1215),
            data_re_in(19) => data_re_in(1279),
            data_re_in(20) => data_re_in(1343),
            data_re_in(21) => data_re_in(1407),
            data_re_in(22) => data_re_in(1471),
            data_re_in(23) => data_re_in(1535),
            data_re_in(24) => data_re_in(1599),
            data_re_in(25) => data_re_in(1663),
            data_re_in(26) => data_re_in(1727),
            data_re_in(27) => data_re_in(1791),
            data_re_in(28) => data_re_in(1855),
            data_re_in(29) => data_re_in(1919),
            data_re_in(30) => data_re_in(1983),
            data_re_in(31) => data_re_in(2047),
            data_im_in(0) => data_im_in(63),
            data_im_in(1) => data_im_in(127),
            data_im_in(2) => data_im_in(191),
            data_im_in(3) => data_im_in(255),
            data_im_in(4) => data_im_in(319),
            data_im_in(5) => data_im_in(383),
            data_im_in(6) => data_im_in(447),
            data_im_in(7) => data_im_in(511),
            data_im_in(8) => data_im_in(575),
            data_im_in(9) => data_im_in(639),
            data_im_in(10) => data_im_in(703),
            data_im_in(11) => data_im_in(767),
            data_im_in(12) => data_im_in(831),
            data_im_in(13) => data_im_in(895),
            data_im_in(14) => data_im_in(959),
            data_im_in(15) => data_im_in(1023),
            data_im_in(16) => data_im_in(1087),
            data_im_in(17) => data_im_in(1151),
            data_im_in(18) => data_im_in(1215),
            data_im_in(19) => data_im_in(1279),
            data_im_in(20) => data_im_in(1343),
            data_im_in(21) => data_im_in(1407),
            data_im_in(22) => data_im_in(1471),
            data_im_in(23) => data_im_in(1535),
            data_im_in(24) => data_im_in(1599),
            data_im_in(25) => data_im_in(1663),
            data_im_in(26) => data_im_in(1727),
            data_im_in(27) => data_im_in(1791),
            data_im_in(28) => data_im_in(1855),
            data_im_in(29) => data_im_in(1919),
            data_im_in(30) => data_im_in(1983),
            data_im_in(31) => data_im_in(2047),
            data_re_out(0) => first_stage_re_out(63),
            data_re_out(1) => first_stage_re_out(127),
            data_re_out(2) => first_stage_re_out(191),
            data_re_out(3) => first_stage_re_out(255),
            data_re_out(4) => first_stage_re_out(319),
            data_re_out(5) => first_stage_re_out(383),
            data_re_out(6) => first_stage_re_out(447),
            data_re_out(7) => first_stage_re_out(511),
            data_re_out(8) => first_stage_re_out(575),
            data_re_out(9) => first_stage_re_out(639),
            data_re_out(10) => first_stage_re_out(703),
            data_re_out(11) => first_stage_re_out(767),
            data_re_out(12) => first_stage_re_out(831),
            data_re_out(13) => first_stage_re_out(895),
            data_re_out(14) => first_stage_re_out(959),
            data_re_out(15) => first_stage_re_out(1023),
            data_re_out(16) => first_stage_re_out(1087),
            data_re_out(17) => first_stage_re_out(1151),
            data_re_out(18) => first_stage_re_out(1215),
            data_re_out(19) => first_stage_re_out(1279),
            data_re_out(20) => first_stage_re_out(1343),
            data_re_out(21) => first_stage_re_out(1407),
            data_re_out(22) => first_stage_re_out(1471),
            data_re_out(23) => first_stage_re_out(1535),
            data_re_out(24) => first_stage_re_out(1599),
            data_re_out(25) => first_stage_re_out(1663),
            data_re_out(26) => first_stage_re_out(1727),
            data_re_out(27) => first_stage_re_out(1791),
            data_re_out(28) => first_stage_re_out(1855),
            data_re_out(29) => first_stage_re_out(1919),
            data_re_out(30) => first_stage_re_out(1983),
            data_re_out(31) => first_stage_re_out(2047),
            data_im_out(0) => first_stage_im_out(63),
            data_im_out(1) => first_stage_im_out(127),
            data_im_out(2) => first_stage_im_out(191),
            data_im_out(3) => first_stage_im_out(255),
            data_im_out(4) => first_stage_im_out(319),
            data_im_out(5) => first_stage_im_out(383),
            data_im_out(6) => first_stage_im_out(447),
            data_im_out(7) => first_stage_im_out(511),
            data_im_out(8) => first_stage_im_out(575),
            data_im_out(9) => first_stage_im_out(639),
            data_im_out(10) => first_stage_im_out(703),
            data_im_out(11) => first_stage_im_out(767),
            data_im_out(12) => first_stage_im_out(831),
            data_im_out(13) => first_stage_im_out(895),
            data_im_out(14) => first_stage_im_out(959),
            data_im_out(15) => first_stage_im_out(1023),
            data_im_out(16) => first_stage_im_out(1087),
            data_im_out(17) => first_stage_im_out(1151),
            data_im_out(18) => first_stage_im_out(1215),
            data_im_out(19) => first_stage_im_out(1279),
            data_im_out(20) => first_stage_im_out(1343),
            data_im_out(21) => first_stage_im_out(1407),
            data_im_out(22) => first_stage_im_out(1471),
            data_im_out(23) => first_stage_im_out(1535),
            data_im_out(24) => first_stage_im_out(1599),
            data_im_out(25) => first_stage_im_out(1663),
            data_im_out(26) => first_stage_im_out(1727),
            data_im_out(27) => first_stage_im_out(1791),
            data_im_out(28) => first_stage_im_out(1855),
            data_im_out(29) => first_stage_im_out(1919),
            data_im_out(30) => first_stage_im_out(1983),
            data_im_out(31) => first_stage_im_out(2047)
        );


    --- right-hand-side processors
    URFFT_PT64_0 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(0),
            data_re_in(1) => mul_re_out(1),
            data_re_in(2) => mul_re_out(2),
            data_re_in(3) => mul_re_out(3),
            data_re_in(4) => mul_re_out(4),
            data_re_in(5) => mul_re_out(5),
            data_re_in(6) => mul_re_out(6),
            data_re_in(7) => mul_re_out(7),
            data_re_in(8) => mul_re_out(8),
            data_re_in(9) => mul_re_out(9),
            data_re_in(10) => mul_re_out(10),
            data_re_in(11) => mul_re_out(11),
            data_re_in(12) => mul_re_out(12),
            data_re_in(13) => mul_re_out(13),
            data_re_in(14) => mul_re_out(14),
            data_re_in(15) => mul_re_out(15),
            data_re_in(16) => mul_re_out(16),
            data_re_in(17) => mul_re_out(17),
            data_re_in(18) => mul_re_out(18),
            data_re_in(19) => mul_re_out(19),
            data_re_in(20) => mul_re_out(20),
            data_re_in(21) => mul_re_out(21),
            data_re_in(22) => mul_re_out(22),
            data_re_in(23) => mul_re_out(23),
            data_re_in(24) => mul_re_out(24),
            data_re_in(25) => mul_re_out(25),
            data_re_in(26) => mul_re_out(26),
            data_re_in(27) => mul_re_out(27),
            data_re_in(28) => mul_re_out(28),
            data_re_in(29) => mul_re_out(29),
            data_re_in(30) => mul_re_out(30),
            data_re_in(31) => mul_re_out(31),
            data_re_in(32) => mul_re_out(32),
            data_re_in(33) => mul_re_out(33),
            data_re_in(34) => mul_re_out(34),
            data_re_in(35) => mul_re_out(35),
            data_re_in(36) => mul_re_out(36),
            data_re_in(37) => mul_re_out(37),
            data_re_in(38) => mul_re_out(38),
            data_re_in(39) => mul_re_out(39),
            data_re_in(40) => mul_re_out(40),
            data_re_in(41) => mul_re_out(41),
            data_re_in(42) => mul_re_out(42),
            data_re_in(43) => mul_re_out(43),
            data_re_in(44) => mul_re_out(44),
            data_re_in(45) => mul_re_out(45),
            data_re_in(46) => mul_re_out(46),
            data_re_in(47) => mul_re_out(47),
            data_re_in(48) => mul_re_out(48),
            data_re_in(49) => mul_re_out(49),
            data_re_in(50) => mul_re_out(50),
            data_re_in(51) => mul_re_out(51),
            data_re_in(52) => mul_re_out(52),
            data_re_in(53) => mul_re_out(53),
            data_re_in(54) => mul_re_out(54),
            data_re_in(55) => mul_re_out(55),
            data_re_in(56) => mul_re_out(56),
            data_re_in(57) => mul_re_out(57),
            data_re_in(58) => mul_re_out(58),
            data_re_in(59) => mul_re_out(59),
            data_re_in(60) => mul_re_out(60),
            data_re_in(61) => mul_re_out(61),
            data_re_in(62) => mul_re_out(62),
            data_re_in(63) => mul_re_out(63),
            data_im_in(0) => mul_im_out(0),
            data_im_in(1) => mul_im_out(1),
            data_im_in(2) => mul_im_out(2),
            data_im_in(3) => mul_im_out(3),
            data_im_in(4) => mul_im_out(4),
            data_im_in(5) => mul_im_out(5),
            data_im_in(6) => mul_im_out(6),
            data_im_in(7) => mul_im_out(7),
            data_im_in(8) => mul_im_out(8),
            data_im_in(9) => mul_im_out(9),
            data_im_in(10) => mul_im_out(10),
            data_im_in(11) => mul_im_out(11),
            data_im_in(12) => mul_im_out(12),
            data_im_in(13) => mul_im_out(13),
            data_im_in(14) => mul_im_out(14),
            data_im_in(15) => mul_im_out(15),
            data_im_in(16) => mul_im_out(16),
            data_im_in(17) => mul_im_out(17),
            data_im_in(18) => mul_im_out(18),
            data_im_in(19) => mul_im_out(19),
            data_im_in(20) => mul_im_out(20),
            data_im_in(21) => mul_im_out(21),
            data_im_in(22) => mul_im_out(22),
            data_im_in(23) => mul_im_out(23),
            data_im_in(24) => mul_im_out(24),
            data_im_in(25) => mul_im_out(25),
            data_im_in(26) => mul_im_out(26),
            data_im_in(27) => mul_im_out(27),
            data_im_in(28) => mul_im_out(28),
            data_im_in(29) => mul_im_out(29),
            data_im_in(30) => mul_im_out(30),
            data_im_in(31) => mul_im_out(31),
            data_im_in(32) => mul_im_out(32),
            data_im_in(33) => mul_im_out(33),
            data_im_in(34) => mul_im_out(34),
            data_im_in(35) => mul_im_out(35),
            data_im_in(36) => mul_im_out(36),
            data_im_in(37) => mul_im_out(37),
            data_im_in(38) => mul_im_out(38),
            data_im_in(39) => mul_im_out(39),
            data_im_in(40) => mul_im_out(40),
            data_im_in(41) => mul_im_out(41),
            data_im_in(42) => mul_im_out(42),
            data_im_in(43) => mul_im_out(43),
            data_im_in(44) => mul_im_out(44),
            data_im_in(45) => mul_im_out(45),
            data_im_in(46) => mul_im_out(46),
            data_im_in(47) => mul_im_out(47),
            data_im_in(48) => mul_im_out(48),
            data_im_in(49) => mul_im_out(49),
            data_im_in(50) => mul_im_out(50),
            data_im_in(51) => mul_im_out(51),
            data_im_in(52) => mul_im_out(52),
            data_im_in(53) => mul_im_out(53),
            data_im_in(54) => mul_im_out(54),
            data_im_in(55) => mul_im_out(55),
            data_im_in(56) => mul_im_out(56),
            data_im_in(57) => mul_im_out(57),
            data_im_in(58) => mul_im_out(58),
            data_im_in(59) => mul_im_out(59),
            data_im_in(60) => mul_im_out(60),
            data_im_in(61) => mul_im_out(61),
            data_im_in(62) => mul_im_out(62),
            data_im_in(63) => mul_im_out(63),
            data_re_out(0) => data_re_out(0),
            data_re_out(1) => data_re_out(32),
            data_re_out(2) => data_re_out(64),
            data_re_out(3) => data_re_out(96),
            data_re_out(4) => data_re_out(128),
            data_re_out(5) => data_re_out(160),
            data_re_out(6) => data_re_out(192),
            data_re_out(7) => data_re_out(224),
            data_re_out(8) => data_re_out(256),
            data_re_out(9) => data_re_out(288),
            data_re_out(10) => data_re_out(320),
            data_re_out(11) => data_re_out(352),
            data_re_out(12) => data_re_out(384),
            data_re_out(13) => data_re_out(416),
            data_re_out(14) => data_re_out(448),
            data_re_out(15) => data_re_out(480),
            data_re_out(16) => data_re_out(512),
            data_re_out(17) => data_re_out(544),
            data_re_out(18) => data_re_out(576),
            data_re_out(19) => data_re_out(608),
            data_re_out(20) => data_re_out(640),
            data_re_out(21) => data_re_out(672),
            data_re_out(22) => data_re_out(704),
            data_re_out(23) => data_re_out(736),
            data_re_out(24) => data_re_out(768),
            data_re_out(25) => data_re_out(800),
            data_re_out(26) => data_re_out(832),
            data_re_out(27) => data_re_out(864),
            data_re_out(28) => data_re_out(896),
            data_re_out(29) => data_re_out(928),
            data_re_out(30) => data_re_out(960),
            data_re_out(31) => data_re_out(992),
            data_re_out(32) => data_re_out(1024),
            data_re_out(33) => data_re_out(1056),
            data_re_out(34) => data_re_out(1088),
            data_re_out(35) => data_re_out(1120),
            data_re_out(36) => data_re_out(1152),
            data_re_out(37) => data_re_out(1184),
            data_re_out(38) => data_re_out(1216),
            data_re_out(39) => data_re_out(1248),
            data_re_out(40) => data_re_out(1280),
            data_re_out(41) => data_re_out(1312),
            data_re_out(42) => data_re_out(1344),
            data_re_out(43) => data_re_out(1376),
            data_re_out(44) => data_re_out(1408),
            data_re_out(45) => data_re_out(1440),
            data_re_out(46) => data_re_out(1472),
            data_re_out(47) => data_re_out(1504),
            data_re_out(48) => data_re_out(1536),
            data_re_out(49) => data_re_out(1568),
            data_re_out(50) => data_re_out(1600),
            data_re_out(51) => data_re_out(1632),
            data_re_out(52) => data_re_out(1664),
            data_re_out(53) => data_re_out(1696),
            data_re_out(54) => data_re_out(1728),
            data_re_out(55) => data_re_out(1760),
            data_re_out(56) => data_re_out(1792),
            data_re_out(57) => data_re_out(1824),
            data_re_out(58) => data_re_out(1856),
            data_re_out(59) => data_re_out(1888),
            data_re_out(60) => data_re_out(1920),
            data_re_out(61) => data_re_out(1952),
            data_re_out(62) => data_re_out(1984),
            data_re_out(63) => data_re_out(2016),
            data_im_out(0) => data_im_out(0),
            data_im_out(1) => data_im_out(32),
            data_im_out(2) => data_im_out(64),
            data_im_out(3) => data_im_out(96),
            data_im_out(4) => data_im_out(128),
            data_im_out(5) => data_im_out(160),
            data_im_out(6) => data_im_out(192),
            data_im_out(7) => data_im_out(224),
            data_im_out(8) => data_im_out(256),
            data_im_out(9) => data_im_out(288),
            data_im_out(10) => data_im_out(320),
            data_im_out(11) => data_im_out(352),
            data_im_out(12) => data_im_out(384),
            data_im_out(13) => data_im_out(416),
            data_im_out(14) => data_im_out(448),
            data_im_out(15) => data_im_out(480),
            data_im_out(16) => data_im_out(512),
            data_im_out(17) => data_im_out(544),
            data_im_out(18) => data_im_out(576),
            data_im_out(19) => data_im_out(608),
            data_im_out(20) => data_im_out(640),
            data_im_out(21) => data_im_out(672),
            data_im_out(22) => data_im_out(704),
            data_im_out(23) => data_im_out(736),
            data_im_out(24) => data_im_out(768),
            data_im_out(25) => data_im_out(800),
            data_im_out(26) => data_im_out(832),
            data_im_out(27) => data_im_out(864),
            data_im_out(28) => data_im_out(896),
            data_im_out(29) => data_im_out(928),
            data_im_out(30) => data_im_out(960),
            data_im_out(31) => data_im_out(992),
            data_im_out(32) => data_im_out(1024),
            data_im_out(33) => data_im_out(1056),
            data_im_out(34) => data_im_out(1088),
            data_im_out(35) => data_im_out(1120),
            data_im_out(36) => data_im_out(1152),
            data_im_out(37) => data_im_out(1184),
            data_im_out(38) => data_im_out(1216),
            data_im_out(39) => data_im_out(1248),
            data_im_out(40) => data_im_out(1280),
            data_im_out(41) => data_im_out(1312),
            data_im_out(42) => data_im_out(1344),
            data_im_out(43) => data_im_out(1376),
            data_im_out(44) => data_im_out(1408),
            data_im_out(45) => data_im_out(1440),
            data_im_out(46) => data_im_out(1472),
            data_im_out(47) => data_im_out(1504),
            data_im_out(48) => data_im_out(1536),
            data_im_out(49) => data_im_out(1568),
            data_im_out(50) => data_im_out(1600),
            data_im_out(51) => data_im_out(1632),
            data_im_out(52) => data_im_out(1664),
            data_im_out(53) => data_im_out(1696),
            data_im_out(54) => data_im_out(1728),
            data_im_out(55) => data_im_out(1760),
            data_im_out(56) => data_im_out(1792),
            data_im_out(57) => data_im_out(1824),
            data_im_out(58) => data_im_out(1856),
            data_im_out(59) => data_im_out(1888),
            data_im_out(60) => data_im_out(1920),
            data_im_out(61) => data_im_out(1952),
            data_im_out(62) => data_im_out(1984),
            data_im_out(63) => data_im_out(2016)
        );           

    URFFT_PT64_1 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(64),
            data_re_in(1) => mul_re_out(65),
            data_re_in(2) => mul_re_out(66),
            data_re_in(3) => mul_re_out(67),
            data_re_in(4) => mul_re_out(68),
            data_re_in(5) => mul_re_out(69),
            data_re_in(6) => mul_re_out(70),
            data_re_in(7) => mul_re_out(71),
            data_re_in(8) => mul_re_out(72),
            data_re_in(9) => mul_re_out(73),
            data_re_in(10) => mul_re_out(74),
            data_re_in(11) => mul_re_out(75),
            data_re_in(12) => mul_re_out(76),
            data_re_in(13) => mul_re_out(77),
            data_re_in(14) => mul_re_out(78),
            data_re_in(15) => mul_re_out(79),
            data_re_in(16) => mul_re_out(80),
            data_re_in(17) => mul_re_out(81),
            data_re_in(18) => mul_re_out(82),
            data_re_in(19) => mul_re_out(83),
            data_re_in(20) => mul_re_out(84),
            data_re_in(21) => mul_re_out(85),
            data_re_in(22) => mul_re_out(86),
            data_re_in(23) => mul_re_out(87),
            data_re_in(24) => mul_re_out(88),
            data_re_in(25) => mul_re_out(89),
            data_re_in(26) => mul_re_out(90),
            data_re_in(27) => mul_re_out(91),
            data_re_in(28) => mul_re_out(92),
            data_re_in(29) => mul_re_out(93),
            data_re_in(30) => mul_re_out(94),
            data_re_in(31) => mul_re_out(95),
            data_re_in(32) => mul_re_out(96),
            data_re_in(33) => mul_re_out(97),
            data_re_in(34) => mul_re_out(98),
            data_re_in(35) => mul_re_out(99),
            data_re_in(36) => mul_re_out(100),
            data_re_in(37) => mul_re_out(101),
            data_re_in(38) => mul_re_out(102),
            data_re_in(39) => mul_re_out(103),
            data_re_in(40) => mul_re_out(104),
            data_re_in(41) => mul_re_out(105),
            data_re_in(42) => mul_re_out(106),
            data_re_in(43) => mul_re_out(107),
            data_re_in(44) => mul_re_out(108),
            data_re_in(45) => mul_re_out(109),
            data_re_in(46) => mul_re_out(110),
            data_re_in(47) => mul_re_out(111),
            data_re_in(48) => mul_re_out(112),
            data_re_in(49) => mul_re_out(113),
            data_re_in(50) => mul_re_out(114),
            data_re_in(51) => mul_re_out(115),
            data_re_in(52) => mul_re_out(116),
            data_re_in(53) => mul_re_out(117),
            data_re_in(54) => mul_re_out(118),
            data_re_in(55) => mul_re_out(119),
            data_re_in(56) => mul_re_out(120),
            data_re_in(57) => mul_re_out(121),
            data_re_in(58) => mul_re_out(122),
            data_re_in(59) => mul_re_out(123),
            data_re_in(60) => mul_re_out(124),
            data_re_in(61) => mul_re_out(125),
            data_re_in(62) => mul_re_out(126),
            data_re_in(63) => mul_re_out(127),
            data_im_in(0) => mul_im_out(64),
            data_im_in(1) => mul_im_out(65),
            data_im_in(2) => mul_im_out(66),
            data_im_in(3) => mul_im_out(67),
            data_im_in(4) => mul_im_out(68),
            data_im_in(5) => mul_im_out(69),
            data_im_in(6) => mul_im_out(70),
            data_im_in(7) => mul_im_out(71),
            data_im_in(8) => mul_im_out(72),
            data_im_in(9) => mul_im_out(73),
            data_im_in(10) => mul_im_out(74),
            data_im_in(11) => mul_im_out(75),
            data_im_in(12) => mul_im_out(76),
            data_im_in(13) => mul_im_out(77),
            data_im_in(14) => mul_im_out(78),
            data_im_in(15) => mul_im_out(79),
            data_im_in(16) => mul_im_out(80),
            data_im_in(17) => mul_im_out(81),
            data_im_in(18) => mul_im_out(82),
            data_im_in(19) => mul_im_out(83),
            data_im_in(20) => mul_im_out(84),
            data_im_in(21) => mul_im_out(85),
            data_im_in(22) => mul_im_out(86),
            data_im_in(23) => mul_im_out(87),
            data_im_in(24) => mul_im_out(88),
            data_im_in(25) => mul_im_out(89),
            data_im_in(26) => mul_im_out(90),
            data_im_in(27) => mul_im_out(91),
            data_im_in(28) => mul_im_out(92),
            data_im_in(29) => mul_im_out(93),
            data_im_in(30) => mul_im_out(94),
            data_im_in(31) => mul_im_out(95),
            data_im_in(32) => mul_im_out(96),
            data_im_in(33) => mul_im_out(97),
            data_im_in(34) => mul_im_out(98),
            data_im_in(35) => mul_im_out(99),
            data_im_in(36) => mul_im_out(100),
            data_im_in(37) => mul_im_out(101),
            data_im_in(38) => mul_im_out(102),
            data_im_in(39) => mul_im_out(103),
            data_im_in(40) => mul_im_out(104),
            data_im_in(41) => mul_im_out(105),
            data_im_in(42) => mul_im_out(106),
            data_im_in(43) => mul_im_out(107),
            data_im_in(44) => mul_im_out(108),
            data_im_in(45) => mul_im_out(109),
            data_im_in(46) => mul_im_out(110),
            data_im_in(47) => mul_im_out(111),
            data_im_in(48) => mul_im_out(112),
            data_im_in(49) => mul_im_out(113),
            data_im_in(50) => mul_im_out(114),
            data_im_in(51) => mul_im_out(115),
            data_im_in(52) => mul_im_out(116),
            data_im_in(53) => mul_im_out(117),
            data_im_in(54) => mul_im_out(118),
            data_im_in(55) => mul_im_out(119),
            data_im_in(56) => mul_im_out(120),
            data_im_in(57) => mul_im_out(121),
            data_im_in(58) => mul_im_out(122),
            data_im_in(59) => mul_im_out(123),
            data_im_in(60) => mul_im_out(124),
            data_im_in(61) => mul_im_out(125),
            data_im_in(62) => mul_im_out(126),
            data_im_in(63) => mul_im_out(127),
            data_re_out(0) => data_re_out(1),
            data_re_out(1) => data_re_out(33),
            data_re_out(2) => data_re_out(65),
            data_re_out(3) => data_re_out(97),
            data_re_out(4) => data_re_out(129),
            data_re_out(5) => data_re_out(161),
            data_re_out(6) => data_re_out(193),
            data_re_out(7) => data_re_out(225),
            data_re_out(8) => data_re_out(257),
            data_re_out(9) => data_re_out(289),
            data_re_out(10) => data_re_out(321),
            data_re_out(11) => data_re_out(353),
            data_re_out(12) => data_re_out(385),
            data_re_out(13) => data_re_out(417),
            data_re_out(14) => data_re_out(449),
            data_re_out(15) => data_re_out(481),
            data_re_out(16) => data_re_out(513),
            data_re_out(17) => data_re_out(545),
            data_re_out(18) => data_re_out(577),
            data_re_out(19) => data_re_out(609),
            data_re_out(20) => data_re_out(641),
            data_re_out(21) => data_re_out(673),
            data_re_out(22) => data_re_out(705),
            data_re_out(23) => data_re_out(737),
            data_re_out(24) => data_re_out(769),
            data_re_out(25) => data_re_out(801),
            data_re_out(26) => data_re_out(833),
            data_re_out(27) => data_re_out(865),
            data_re_out(28) => data_re_out(897),
            data_re_out(29) => data_re_out(929),
            data_re_out(30) => data_re_out(961),
            data_re_out(31) => data_re_out(993),
            data_re_out(32) => data_re_out(1025),
            data_re_out(33) => data_re_out(1057),
            data_re_out(34) => data_re_out(1089),
            data_re_out(35) => data_re_out(1121),
            data_re_out(36) => data_re_out(1153),
            data_re_out(37) => data_re_out(1185),
            data_re_out(38) => data_re_out(1217),
            data_re_out(39) => data_re_out(1249),
            data_re_out(40) => data_re_out(1281),
            data_re_out(41) => data_re_out(1313),
            data_re_out(42) => data_re_out(1345),
            data_re_out(43) => data_re_out(1377),
            data_re_out(44) => data_re_out(1409),
            data_re_out(45) => data_re_out(1441),
            data_re_out(46) => data_re_out(1473),
            data_re_out(47) => data_re_out(1505),
            data_re_out(48) => data_re_out(1537),
            data_re_out(49) => data_re_out(1569),
            data_re_out(50) => data_re_out(1601),
            data_re_out(51) => data_re_out(1633),
            data_re_out(52) => data_re_out(1665),
            data_re_out(53) => data_re_out(1697),
            data_re_out(54) => data_re_out(1729),
            data_re_out(55) => data_re_out(1761),
            data_re_out(56) => data_re_out(1793),
            data_re_out(57) => data_re_out(1825),
            data_re_out(58) => data_re_out(1857),
            data_re_out(59) => data_re_out(1889),
            data_re_out(60) => data_re_out(1921),
            data_re_out(61) => data_re_out(1953),
            data_re_out(62) => data_re_out(1985),
            data_re_out(63) => data_re_out(2017),
            data_im_out(0) => data_im_out(1),
            data_im_out(1) => data_im_out(33),
            data_im_out(2) => data_im_out(65),
            data_im_out(3) => data_im_out(97),
            data_im_out(4) => data_im_out(129),
            data_im_out(5) => data_im_out(161),
            data_im_out(6) => data_im_out(193),
            data_im_out(7) => data_im_out(225),
            data_im_out(8) => data_im_out(257),
            data_im_out(9) => data_im_out(289),
            data_im_out(10) => data_im_out(321),
            data_im_out(11) => data_im_out(353),
            data_im_out(12) => data_im_out(385),
            data_im_out(13) => data_im_out(417),
            data_im_out(14) => data_im_out(449),
            data_im_out(15) => data_im_out(481),
            data_im_out(16) => data_im_out(513),
            data_im_out(17) => data_im_out(545),
            data_im_out(18) => data_im_out(577),
            data_im_out(19) => data_im_out(609),
            data_im_out(20) => data_im_out(641),
            data_im_out(21) => data_im_out(673),
            data_im_out(22) => data_im_out(705),
            data_im_out(23) => data_im_out(737),
            data_im_out(24) => data_im_out(769),
            data_im_out(25) => data_im_out(801),
            data_im_out(26) => data_im_out(833),
            data_im_out(27) => data_im_out(865),
            data_im_out(28) => data_im_out(897),
            data_im_out(29) => data_im_out(929),
            data_im_out(30) => data_im_out(961),
            data_im_out(31) => data_im_out(993),
            data_im_out(32) => data_im_out(1025),
            data_im_out(33) => data_im_out(1057),
            data_im_out(34) => data_im_out(1089),
            data_im_out(35) => data_im_out(1121),
            data_im_out(36) => data_im_out(1153),
            data_im_out(37) => data_im_out(1185),
            data_im_out(38) => data_im_out(1217),
            data_im_out(39) => data_im_out(1249),
            data_im_out(40) => data_im_out(1281),
            data_im_out(41) => data_im_out(1313),
            data_im_out(42) => data_im_out(1345),
            data_im_out(43) => data_im_out(1377),
            data_im_out(44) => data_im_out(1409),
            data_im_out(45) => data_im_out(1441),
            data_im_out(46) => data_im_out(1473),
            data_im_out(47) => data_im_out(1505),
            data_im_out(48) => data_im_out(1537),
            data_im_out(49) => data_im_out(1569),
            data_im_out(50) => data_im_out(1601),
            data_im_out(51) => data_im_out(1633),
            data_im_out(52) => data_im_out(1665),
            data_im_out(53) => data_im_out(1697),
            data_im_out(54) => data_im_out(1729),
            data_im_out(55) => data_im_out(1761),
            data_im_out(56) => data_im_out(1793),
            data_im_out(57) => data_im_out(1825),
            data_im_out(58) => data_im_out(1857),
            data_im_out(59) => data_im_out(1889),
            data_im_out(60) => data_im_out(1921),
            data_im_out(61) => data_im_out(1953),
            data_im_out(62) => data_im_out(1985),
            data_im_out(63) => data_im_out(2017)
        );           

    URFFT_PT64_2 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(128),
            data_re_in(1) => mul_re_out(129),
            data_re_in(2) => mul_re_out(130),
            data_re_in(3) => mul_re_out(131),
            data_re_in(4) => mul_re_out(132),
            data_re_in(5) => mul_re_out(133),
            data_re_in(6) => mul_re_out(134),
            data_re_in(7) => mul_re_out(135),
            data_re_in(8) => mul_re_out(136),
            data_re_in(9) => mul_re_out(137),
            data_re_in(10) => mul_re_out(138),
            data_re_in(11) => mul_re_out(139),
            data_re_in(12) => mul_re_out(140),
            data_re_in(13) => mul_re_out(141),
            data_re_in(14) => mul_re_out(142),
            data_re_in(15) => mul_re_out(143),
            data_re_in(16) => mul_re_out(144),
            data_re_in(17) => mul_re_out(145),
            data_re_in(18) => mul_re_out(146),
            data_re_in(19) => mul_re_out(147),
            data_re_in(20) => mul_re_out(148),
            data_re_in(21) => mul_re_out(149),
            data_re_in(22) => mul_re_out(150),
            data_re_in(23) => mul_re_out(151),
            data_re_in(24) => mul_re_out(152),
            data_re_in(25) => mul_re_out(153),
            data_re_in(26) => mul_re_out(154),
            data_re_in(27) => mul_re_out(155),
            data_re_in(28) => mul_re_out(156),
            data_re_in(29) => mul_re_out(157),
            data_re_in(30) => mul_re_out(158),
            data_re_in(31) => mul_re_out(159),
            data_re_in(32) => mul_re_out(160),
            data_re_in(33) => mul_re_out(161),
            data_re_in(34) => mul_re_out(162),
            data_re_in(35) => mul_re_out(163),
            data_re_in(36) => mul_re_out(164),
            data_re_in(37) => mul_re_out(165),
            data_re_in(38) => mul_re_out(166),
            data_re_in(39) => mul_re_out(167),
            data_re_in(40) => mul_re_out(168),
            data_re_in(41) => mul_re_out(169),
            data_re_in(42) => mul_re_out(170),
            data_re_in(43) => mul_re_out(171),
            data_re_in(44) => mul_re_out(172),
            data_re_in(45) => mul_re_out(173),
            data_re_in(46) => mul_re_out(174),
            data_re_in(47) => mul_re_out(175),
            data_re_in(48) => mul_re_out(176),
            data_re_in(49) => mul_re_out(177),
            data_re_in(50) => mul_re_out(178),
            data_re_in(51) => mul_re_out(179),
            data_re_in(52) => mul_re_out(180),
            data_re_in(53) => mul_re_out(181),
            data_re_in(54) => mul_re_out(182),
            data_re_in(55) => mul_re_out(183),
            data_re_in(56) => mul_re_out(184),
            data_re_in(57) => mul_re_out(185),
            data_re_in(58) => mul_re_out(186),
            data_re_in(59) => mul_re_out(187),
            data_re_in(60) => mul_re_out(188),
            data_re_in(61) => mul_re_out(189),
            data_re_in(62) => mul_re_out(190),
            data_re_in(63) => mul_re_out(191),
            data_im_in(0) => mul_im_out(128),
            data_im_in(1) => mul_im_out(129),
            data_im_in(2) => mul_im_out(130),
            data_im_in(3) => mul_im_out(131),
            data_im_in(4) => mul_im_out(132),
            data_im_in(5) => mul_im_out(133),
            data_im_in(6) => mul_im_out(134),
            data_im_in(7) => mul_im_out(135),
            data_im_in(8) => mul_im_out(136),
            data_im_in(9) => mul_im_out(137),
            data_im_in(10) => mul_im_out(138),
            data_im_in(11) => mul_im_out(139),
            data_im_in(12) => mul_im_out(140),
            data_im_in(13) => mul_im_out(141),
            data_im_in(14) => mul_im_out(142),
            data_im_in(15) => mul_im_out(143),
            data_im_in(16) => mul_im_out(144),
            data_im_in(17) => mul_im_out(145),
            data_im_in(18) => mul_im_out(146),
            data_im_in(19) => mul_im_out(147),
            data_im_in(20) => mul_im_out(148),
            data_im_in(21) => mul_im_out(149),
            data_im_in(22) => mul_im_out(150),
            data_im_in(23) => mul_im_out(151),
            data_im_in(24) => mul_im_out(152),
            data_im_in(25) => mul_im_out(153),
            data_im_in(26) => mul_im_out(154),
            data_im_in(27) => mul_im_out(155),
            data_im_in(28) => mul_im_out(156),
            data_im_in(29) => mul_im_out(157),
            data_im_in(30) => mul_im_out(158),
            data_im_in(31) => mul_im_out(159),
            data_im_in(32) => mul_im_out(160),
            data_im_in(33) => mul_im_out(161),
            data_im_in(34) => mul_im_out(162),
            data_im_in(35) => mul_im_out(163),
            data_im_in(36) => mul_im_out(164),
            data_im_in(37) => mul_im_out(165),
            data_im_in(38) => mul_im_out(166),
            data_im_in(39) => mul_im_out(167),
            data_im_in(40) => mul_im_out(168),
            data_im_in(41) => mul_im_out(169),
            data_im_in(42) => mul_im_out(170),
            data_im_in(43) => mul_im_out(171),
            data_im_in(44) => mul_im_out(172),
            data_im_in(45) => mul_im_out(173),
            data_im_in(46) => mul_im_out(174),
            data_im_in(47) => mul_im_out(175),
            data_im_in(48) => mul_im_out(176),
            data_im_in(49) => mul_im_out(177),
            data_im_in(50) => mul_im_out(178),
            data_im_in(51) => mul_im_out(179),
            data_im_in(52) => mul_im_out(180),
            data_im_in(53) => mul_im_out(181),
            data_im_in(54) => mul_im_out(182),
            data_im_in(55) => mul_im_out(183),
            data_im_in(56) => mul_im_out(184),
            data_im_in(57) => mul_im_out(185),
            data_im_in(58) => mul_im_out(186),
            data_im_in(59) => mul_im_out(187),
            data_im_in(60) => mul_im_out(188),
            data_im_in(61) => mul_im_out(189),
            data_im_in(62) => mul_im_out(190),
            data_im_in(63) => mul_im_out(191),
            data_re_out(0) => data_re_out(2),
            data_re_out(1) => data_re_out(34),
            data_re_out(2) => data_re_out(66),
            data_re_out(3) => data_re_out(98),
            data_re_out(4) => data_re_out(130),
            data_re_out(5) => data_re_out(162),
            data_re_out(6) => data_re_out(194),
            data_re_out(7) => data_re_out(226),
            data_re_out(8) => data_re_out(258),
            data_re_out(9) => data_re_out(290),
            data_re_out(10) => data_re_out(322),
            data_re_out(11) => data_re_out(354),
            data_re_out(12) => data_re_out(386),
            data_re_out(13) => data_re_out(418),
            data_re_out(14) => data_re_out(450),
            data_re_out(15) => data_re_out(482),
            data_re_out(16) => data_re_out(514),
            data_re_out(17) => data_re_out(546),
            data_re_out(18) => data_re_out(578),
            data_re_out(19) => data_re_out(610),
            data_re_out(20) => data_re_out(642),
            data_re_out(21) => data_re_out(674),
            data_re_out(22) => data_re_out(706),
            data_re_out(23) => data_re_out(738),
            data_re_out(24) => data_re_out(770),
            data_re_out(25) => data_re_out(802),
            data_re_out(26) => data_re_out(834),
            data_re_out(27) => data_re_out(866),
            data_re_out(28) => data_re_out(898),
            data_re_out(29) => data_re_out(930),
            data_re_out(30) => data_re_out(962),
            data_re_out(31) => data_re_out(994),
            data_re_out(32) => data_re_out(1026),
            data_re_out(33) => data_re_out(1058),
            data_re_out(34) => data_re_out(1090),
            data_re_out(35) => data_re_out(1122),
            data_re_out(36) => data_re_out(1154),
            data_re_out(37) => data_re_out(1186),
            data_re_out(38) => data_re_out(1218),
            data_re_out(39) => data_re_out(1250),
            data_re_out(40) => data_re_out(1282),
            data_re_out(41) => data_re_out(1314),
            data_re_out(42) => data_re_out(1346),
            data_re_out(43) => data_re_out(1378),
            data_re_out(44) => data_re_out(1410),
            data_re_out(45) => data_re_out(1442),
            data_re_out(46) => data_re_out(1474),
            data_re_out(47) => data_re_out(1506),
            data_re_out(48) => data_re_out(1538),
            data_re_out(49) => data_re_out(1570),
            data_re_out(50) => data_re_out(1602),
            data_re_out(51) => data_re_out(1634),
            data_re_out(52) => data_re_out(1666),
            data_re_out(53) => data_re_out(1698),
            data_re_out(54) => data_re_out(1730),
            data_re_out(55) => data_re_out(1762),
            data_re_out(56) => data_re_out(1794),
            data_re_out(57) => data_re_out(1826),
            data_re_out(58) => data_re_out(1858),
            data_re_out(59) => data_re_out(1890),
            data_re_out(60) => data_re_out(1922),
            data_re_out(61) => data_re_out(1954),
            data_re_out(62) => data_re_out(1986),
            data_re_out(63) => data_re_out(2018),
            data_im_out(0) => data_im_out(2),
            data_im_out(1) => data_im_out(34),
            data_im_out(2) => data_im_out(66),
            data_im_out(3) => data_im_out(98),
            data_im_out(4) => data_im_out(130),
            data_im_out(5) => data_im_out(162),
            data_im_out(6) => data_im_out(194),
            data_im_out(7) => data_im_out(226),
            data_im_out(8) => data_im_out(258),
            data_im_out(9) => data_im_out(290),
            data_im_out(10) => data_im_out(322),
            data_im_out(11) => data_im_out(354),
            data_im_out(12) => data_im_out(386),
            data_im_out(13) => data_im_out(418),
            data_im_out(14) => data_im_out(450),
            data_im_out(15) => data_im_out(482),
            data_im_out(16) => data_im_out(514),
            data_im_out(17) => data_im_out(546),
            data_im_out(18) => data_im_out(578),
            data_im_out(19) => data_im_out(610),
            data_im_out(20) => data_im_out(642),
            data_im_out(21) => data_im_out(674),
            data_im_out(22) => data_im_out(706),
            data_im_out(23) => data_im_out(738),
            data_im_out(24) => data_im_out(770),
            data_im_out(25) => data_im_out(802),
            data_im_out(26) => data_im_out(834),
            data_im_out(27) => data_im_out(866),
            data_im_out(28) => data_im_out(898),
            data_im_out(29) => data_im_out(930),
            data_im_out(30) => data_im_out(962),
            data_im_out(31) => data_im_out(994),
            data_im_out(32) => data_im_out(1026),
            data_im_out(33) => data_im_out(1058),
            data_im_out(34) => data_im_out(1090),
            data_im_out(35) => data_im_out(1122),
            data_im_out(36) => data_im_out(1154),
            data_im_out(37) => data_im_out(1186),
            data_im_out(38) => data_im_out(1218),
            data_im_out(39) => data_im_out(1250),
            data_im_out(40) => data_im_out(1282),
            data_im_out(41) => data_im_out(1314),
            data_im_out(42) => data_im_out(1346),
            data_im_out(43) => data_im_out(1378),
            data_im_out(44) => data_im_out(1410),
            data_im_out(45) => data_im_out(1442),
            data_im_out(46) => data_im_out(1474),
            data_im_out(47) => data_im_out(1506),
            data_im_out(48) => data_im_out(1538),
            data_im_out(49) => data_im_out(1570),
            data_im_out(50) => data_im_out(1602),
            data_im_out(51) => data_im_out(1634),
            data_im_out(52) => data_im_out(1666),
            data_im_out(53) => data_im_out(1698),
            data_im_out(54) => data_im_out(1730),
            data_im_out(55) => data_im_out(1762),
            data_im_out(56) => data_im_out(1794),
            data_im_out(57) => data_im_out(1826),
            data_im_out(58) => data_im_out(1858),
            data_im_out(59) => data_im_out(1890),
            data_im_out(60) => data_im_out(1922),
            data_im_out(61) => data_im_out(1954),
            data_im_out(62) => data_im_out(1986),
            data_im_out(63) => data_im_out(2018)
        );           

    URFFT_PT64_3 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(192),
            data_re_in(1) => mul_re_out(193),
            data_re_in(2) => mul_re_out(194),
            data_re_in(3) => mul_re_out(195),
            data_re_in(4) => mul_re_out(196),
            data_re_in(5) => mul_re_out(197),
            data_re_in(6) => mul_re_out(198),
            data_re_in(7) => mul_re_out(199),
            data_re_in(8) => mul_re_out(200),
            data_re_in(9) => mul_re_out(201),
            data_re_in(10) => mul_re_out(202),
            data_re_in(11) => mul_re_out(203),
            data_re_in(12) => mul_re_out(204),
            data_re_in(13) => mul_re_out(205),
            data_re_in(14) => mul_re_out(206),
            data_re_in(15) => mul_re_out(207),
            data_re_in(16) => mul_re_out(208),
            data_re_in(17) => mul_re_out(209),
            data_re_in(18) => mul_re_out(210),
            data_re_in(19) => mul_re_out(211),
            data_re_in(20) => mul_re_out(212),
            data_re_in(21) => mul_re_out(213),
            data_re_in(22) => mul_re_out(214),
            data_re_in(23) => mul_re_out(215),
            data_re_in(24) => mul_re_out(216),
            data_re_in(25) => mul_re_out(217),
            data_re_in(26) => mul_re_out(218),
            data_re_in(27) => mul_re_out(219),
            data_re_in(28) => mul_re_out(220),
            data_re_in(29) => mul_re_out(221),
            data_re_in(30) => mul_re_out(222),
            data_re_in(31) => mul_re_out(223),
            data_re_in(32) => mul_re_out(224),
            data_re_in(33) => mul_re_out(225),
            data_re_in(34) => mul_re_out(226),
            data_re_in(35) => mul_re_out(227),
            data_re_in(36) => mul_re_out(228),
            data_re_in(37) => mul_re_out(229),
            data_re_in(38) => mul_re_out(230),
            data_re_in(39) => mul_re_out(231),
            data_re_in(40) => mul_re_out(232),
            data_re_in(41) => mul_re_out(233),
            data_re_in(42) => mul_re_out(234),
            data_re_in(43) => mul_re_out(235),
            data_re_in(44) => mul_re_out(236),
            data_re_in(45) => mul_re_out(237),
            data_re_in(46) => mul_re_out(238),
            data_re_in(47) => mul_re_out(239),
            data_re_in(48) => mul_re_out(240),
            data_re_in(49) => mul_re_out(241),
            data_re_in(50) => mul_re_out(242),
            data_re_in(51) => mul_re_out(243),
            data_re_in(52) => mul_re_out(244),
            data_re_in(53) => mul_re_out(245),
            data_re_in(54) => mul_re_out(246),
            data_re_in(55) => mul_re_out(247),
            data_re_in(56) => mul_re_out(248),
            data_re_in(57) => mul_re_out(249),
            data_re_in(58) => mul_re_out(250),
            data_re_in(59) => mul_re_out(251),
            data_re_in(60) => mul_re_out(252),
            data_re_in(61) => mul_re_out(253),
            data_re_in(62) => mul_re_out(254),
            data_re_in(63) => mul_re_out(255),
            data_im_in(0) => mul_im_out(192),
            data_im_in(1) => mul_im_out(193),
            data_im_in(2) => mul_im_out(194),
            data_im_in(3) => mul_im_out(195),
            data_im_in(4) => mul_im_out(196),
            data_im_in(5) => mul_im_out(197),
            data_im_in(6) => mul_im_out(198),
            data_im_in(7) => mul_im_out(199),
            data_im_in(8) => mul_im_out(200),
            data_im_in(9) => mul_im_out(201),
            data_im_in(10) => mul_im_out(202),
            data_im_in(11) => mul_im_out(203),
            data_im_in(12) => mul_im_out(204),
            data_im_in(13) => mul_im_out(205),
            data_im_in(14) => mul_im_out(206),
            data_im_in(15) => mul_im_out(207),
            data_im_in(16) => mul_im_out(208),
            data_im_in(17) => mul_im_out(209),
            data_im_in(18) => mul_im_out(210),
            data_im_in(19) => mul_im_out(211),
            data_im_in(20) => mul_im_out(212),
            data_im_in(21) => mul_im_out(213),
            data_im_in(22) => mul_im_out(214),
            data_im_in(23) => mul_im_out(215),
            data_im_in(24) => mul_im_out(216),
            data_im_in(25) => mul_im_out(217),
            data_im_in(26) => mul_im_out(218),
            data_im_in(27) => mul_im_out(219),
            data_im_in(28) => mul_im_out(220),
            data_im_in(29) => mul_im_out(221),
            data_im_in(30) => mul_im_out(222),
            data_im_in(31) => mul_im_out(223),
            data_im_in(32) => mul_im_out(224),
            data_im_in(33) => mul_im_out(225),
            data_im_in(34) => mul_im_out(226),
            data_im_in(35) => mul_im_out(227),
            data_im_in(36) => mul_im_out(228),
            data_im_in(37) => mul_im_out(229),
            data_im_in(38) => mul_im_out(230),
            data_im_in(39) => mul_im_out(231),
            data_im_in(40) => mul_im_out(232),
            data_im_in(41) => mul_im_out(233),
            data_im_in(42) => mul_im_out(234),
            data_im_in(43) => mul_im_out(235),
            data_im_in(44) => mul_im_out(236),
            data_im_in(45) => mul_im_out(237),
            data_im_in(46) => mul_im_out(238),
            data_im_in(47) => mul_im_out(239),
            data_im_in(48) => mul_im_out(240),
            data_im_in(49) => mul_im_out(241),
            data_im_in(50) => mul_im_out(242),
            data_im_in(51) => mul_im_out(243),
            data_im_in(52) => mul_im_out(244),
            data_im_in(53) => mul_im_out(245),
            data_im_in(54) => mul_im_out(246),
            data_im_in(55) => mul_im_out(247),
            data_im_in(56) => mul_im_out(248),
            data_im_in(57) => mul_im_out(249),
            data_im_in(58) => mul_im_out(250),
            data_im_in(59) => mul_im_out(251),
            data_im_in(60) => mul_im_out(252),
            data_im_in(61) => mul_im_out(253),
            data_im_in(62) => mul_im_out(254),
            data_im_in(63) => mul_im_out(255),
            data_re_out(0) => data_re_out(3),
            data_re_out(1) => data_re_out(35),
            data_re_out(2) => data_re_out(67),
            data_re_out(3) => data_re_out(99),
            data_re_out(4) => data_re_out(131),
            data_re_out(5) => data_re_out(163),
            data_re_out(6) => data_re_out(195),
            data_re_out(7) => data_re_out(227),
            data_re_out(8) => data_re_out(259),
            data_re_out(9) => data_re_out(291),
            data_re_out(10) => data_re_out(323),
            data_re_out(11) => data_re_out(355),
            data_re_out(12) => data_re_out(387),
            data_re_out(13) => data_re_out(419),
            data_re_out(14) => data_re_out(451),
            data_re_out(15) => data_re_out(483),
            data_re_out(16) => data_re_out(515),
            data_re_out(17) => data_re_out(547),
            data_re_out(18) => data_re_out(579),
            data_re_out(19) => data_re_out(611),
            data_re_out(20) => data_re_out(643),
            data_re_out(21) => data_re_out(675),
            data_re_out(22) => data_re_out(707),
            data_re_out(23) => data_re_out(739),
            data_re_out(24) => data_re_out(771),
            data_re_out(25) => data_re_out(803),
            data_re_out(26) => data_re_out(835),
            data_re_out(27) => data_re_out(867),
            data_re_out(28) => data_re_out(899),
            data_re_out(29) => data_re_out(931),
            data_re_out(30) => data_re_out(963),
            data_re_out(31) => data_re_out(995),
            data_re_out(32) => data_re_out(1027),
            data_re_out(33) => data_re_out(1059),
            data_re_out(34) => data_re_out(1091),
            data_re_out(35) => data_re_out(1123),
            data_re_out(36) => data_re_out(1155),
            data_re_out(37) => data_re_out(1187),
            data_re_out(38) => data_re_out(1219),
            data_re_out(39) => data_re_out(1251),
            data_re_out(40) => data_re_out(1283),
            data_re_out(41) => data_re_out(1315),
            data_re_out(42) => data_re_out(1347),
            data_re_out(43) => data_re_out(1379),
            data_re_out(44) => data_re_out(1411),
            data_re_out(45) => data_re_out(1443),
            data_re_out(46) => data_re_out(1475),
            data_re_out(47) => data_re_out(1507),
            data_re_out(48) => data_re_out(1539),
            data_re_out(49) => data_re_out(1571),
            data_re_out(50) => data_re_out(1603),
            data_re_out(51) => data_re_out(1635),
            data_re_out(52) => data_re_out(1667),
            data_re_out(53) => data_re_out(1699),
            data_re_out(54) => data_re_out(1731),
            data_re_out(55) => data_re_out(1763),
            data_re_out(56) => data_re_out(1795),
            data_re_out(57) => data_re_out(1827),
            data_re_out(58) => data_re_out(1859),
            data_re_out(59) => data_re_out(1891),
            data_re_out(60) => data_re_out(1923),
            data_re_out(61) => data_re_out(1955),
            data_re_out(62) => data_re_out(1987),
            data_re_out(63) => data_re_out(2019),
            data_im_out(0) => data_im_out(3),
            data_im_out(1) => data_im_out(35),
            data_im_out(2) => data_im_out(67),
            data_im_out(3) => data_im_out(99),
            data_im_out(4) => data_im_out(131),
            data_im_out(5) => data_im_out(163),
            data_im_out(6) => data_im_out(195),
            data_im_out(7) => data_im_out(227),
            data_im_out(8) => data_im_out(259),
            data_im_out(9) => data_im_out(291),
            data_im_out(10) => data_im_out(323),
            data_im_out(11) => data_im_out(355),
            data_im_out(12) => data_im_out(387),
            data_im_out(13) => data_im_out(419),
            data_im_out(14) => data_im_out(451),
            data_im_out(15) => data_im_out(483),
            data_im_out(16) => data_im_out(515),
            data_im_out(17) => data_im_out(547),
            data_im_out(18) => data_im_out(579),
            data_im_out(19) => data_im_out(611),
            data_im_out(20) => data_im_out(643),
            data_im_out(21) => data_im_out(675),
            data_im_out(22) => data_im_out(707),
            data_im_out(23) => data_im_out(739),
            data_im_out(24) => data_im_out(771),
            data_im_out(25) => data_im_out(803),
            data_im_out(26) => data_im_out(835),
            data_im_out(27) => data_im_out(867),
            data_im_out(28) => data_im_out(899),
            data_im_out(29) => data_im_out(931),
            data_im_out(30) => data_im_out(963),
            data_im_out(31) => data_im_out(995),
            data_im_out(32) => data_im_out(1027),
            data_im_out(33) => data_im_out(1059),
            data_im_out(34) => data_im_out(1091),
            data_im_out(35) => data_im_out(1123),
            data_im_out(36) => data_im_out(1155),
            data_im_out(37) => data_im_out(1187),
            data_im_out(38) => data_im_out(1219),
            data_im_out(39) => data_im_out(1251),
            data_im_out(40) => data_im_out(1283),
            data_im_out(41) => data_im_out(1315),
            data_im_out(42) => data_im_out(1347),
            data_im_out(43) => data_im_out(1379),
            data_im_out(44) => data_im_out(1411),
            data_im_out(45) => data_im_out(1443),
            data_im_out(46) => data_im_out(1475),
            data_im_out(47) => data_im_out(1507),
            data_im_out(48) => data_im_out(1539),
            data_im_out(49) => data_im_out(1571),
            data_im_out(50) => data_im_out(1603),
            data_im_out(51) => data_im_out(1635),
            data_im_out(52) => data_im_out(1667),
            data_im_out(53) => data_im_out(1699),
            data_im_out(54) => data_im_out(1731),
            data_im_out(55) => data_im_out(1763),
            data_im_out(56) => data_im_out(1795),
            data_im_out(57) => data_im_out(1827),
            data_im_out(58) => data_im_out(1859),
            data_im_out(59) => data_im_out(1891),
            data_im_out(60) => data_im_out(1923),
            data_im_out(61) => data_im_out(1955),
            data_im_out(62) => data_im_out(1987),
            data_im_out(63) => data_im_out(2019)
        );           

    URFFT_PT64_4 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(256),
            data_re_in(1) => mul_re_out(257),
            data_re_in(2) => mul_re_out(258),
            data_re_in(3) => mul_re_out(259),
            data_re_in(4) => mul_re_out(260),
            data_re_in(5) => mul_re_out(261),
            data_re_in(6) => mul_re_out(262),
            data_re_in(7) => mul_re_out(263),
            data_re_in(8) => mul_re_out(264),
            data_re_in(9) => mul_re_out(265),
            data_re_in(10) => mul_re_out(266),
            data_re_in(11) => mul_re_out(267),
            data_re_in(12) => mul_re_out(268),
            data_re_in(13) => mul_re_out(269),
            data_re_in(14) => mul_re_out(270),
            data_re_in(15) => mul_re_out(271),
            data_re_in(16) => mul_re_out(272),
            data_re_in(17) => mul_re_out(273),
            data_re_in(18) => mul_re_out(274),
            data_re_in(19) => mul_re_out(275),
            data_re_in(20) => mul_re_out(276),
            data_re_in(21) => mul_re_out(277),
            data_re_in(22) => mul_re_out(278),
            data_re_in(23) => mul_re_out(279),
            data_re_in(24) => mul_re_out(280),
            data_re_in(25) => mul_re_out(281),
            data_re_in(26) => mul_re_out(282),
            data_re_in(27) => mul_re_out(283),
            data_re_in(28) => mul_re_out(284),
            data_re_in(29) => mul_re_out(285),
            data_re_in(30) => mul_re_out(286),
            data_re_in(31) => mul_re_out(287),
            data_re_in(32) => mul_re_out(288),
            data_re_in(33) => mul_re_out(289),
            data_re_in(34) => mul_re_out(290),
            data_re_in(35) => mul_re_out(291),
            data_re_in(36) => mul_re_out(292),
            data_re_in(37) => mul_re_out(293),
            data_re_in(38) => mul_re_out(294),
            data_re_in(39) => mul_re_out(295),
            data_re_in(40) => mul_re_out(296),
            data_re_in(41) => mul_re_out(297),
            data_re_in(42) => mul_re_out(298),
            data_re_in(43) => mul_re_out(299),
            data_re_in(44) => mul_re_out(300),
            data_re_in(45) => mul_re_out(301),
            data_re_in(46) => mul_re_out(302),
            data_re_in(47) => mul_re_out(303),
            data_re_in(48) => mul_re_out(304),
            data_re_in(49) => mul_re_out(305),
            data_re_in(50) => mul_re_out(306),
            data_re_in(51) => mul_re_out(307),
            data_re_in(52) => mul_re_out(308),
            data_re_in(53) => mul_re_out(309),
            data_re_in(54) => mul_re_out(310),
            data_re_in(55) => mul_re_out(311),
            data_re_in(56) => mul_re_out(312),
            data_re_in(57) => mul_re_out(313),
            data_re_in(58) => mul_re_out(314),
            data_re_in(59) => mul_re_out(315),
            data_re_in(60) => mul_re_out(316),
            data_re_in(61) => mul_re_out(317),
            data_re_in(62) => mul_re_out(318),
            data_re_in(63) => mul_re_out(319),
            data_im_in(0) => mul_im_out(256),
            data_im_in(1) => mul_im_out(257),
            data_im_in(2) => mul_im_out(258),
            data_im_in(3) => mul_im_out(259),
            data_im_in(4) => mul_im_out(260),
            data_im_in(5) => mul_im_out(261),
            data_im_in(6) => mul_im_out(262),
            data_im_in(7) => mul_im_out(263),
            data_im_in(8) => mul_im_out(264),
            data_im_in(9) => mul_im_out(265),
            data_im_in(10) => mul_im_out(266),
            data_im_in(11) => mul_im_out(267),
            data_im_in(12) => mul_im_out(268),
            data_im_in(13) => mul_im_out(269),
            data_im_in(14) => mul_im_out(270),
            data_im_in(15) => mul_im_out(271),
            data_im_in(16) => mul_im_out(272),
            data_im_in(17) => mul_im_out(273),
            data_im_in(18) => mul_im_out(274),
            data_im_in(19) => mul_im_out(275),
            data_im_in(20) => mul_im_out(276),
            data_im_in(21) => mul_im_out(277),
            data_im_in(22) => mul_im_out(278),
            data_im_in(23) => mul_im_out(279),
            data_im_in(24) => mul_im_out(280),
            data_im_in(25) => mul_im_out(281),
            data_im_in(26) => mul_im_out(282),
            data_im_in(27) => mul_im_out(283),
            data_im_in(28) => mul_im_out(284),
            data_im_in(29) => mul_im_out(285),
            data_im_in(30) => mul_im_out(286),
            data_im_in(31) => mul_im_out(287),
            data_im_in(32) => mul_im_out(288),
            data_im_in(33) => mul_im_out(289),
            data_im_in(34) => mul_im_out(290),
            data_im_in(35) => mul_im_out(291),
            data_im_in(36) => mul_im_out(292),
            data_im_in(37) => mul_im_out(293),
            data_im_in(38) => mul_im_out(294),
            data_im_in(39) => mul_im_out(295),
            data_im_in(40) => mul_im_out(296),
            data_im_in(41) => mul_im_out(297),
            data_im_in(42) => mul_im_out(298),
            data_im_in(43) => mul_im_out(299),
            data_im_in(44) => mul_im_out(300),
            data_im_in(45) => mul_im_out(301),
            data_im_in(46) => mul_im_out(302),
            data_im_in(47) => mul_im_out(303),
            data_im_in(48) => mul_im_out(304),
            data_im_in(49) => mul_im_out(305),
            data_im_in(50) => mul_im_out(306),
            data_im_in(51) => mul_im_out(307),
            data_im_in(52) => mul_im_out(308),
            data_im_in(53) => mul_im_out(309),
            data_im_in(54) => mul_im_out(310),
            data_im_in(55) => mul_im_out(311),
            data_im_in(56) => mul_im_out(312),
            data_im_in(57) => mul_im_out(313),
            data_im_in(58) => mul_im_out(314),
            data_im_in(59) => mul_im_out(315),
            data_im_in(60) => mul_im_out(316),
            data_im_in(61) => mul_im_out(317),
            data_im_in(62) => mul_im_out(318),
            data_im_in(63) => mul_im_out(319),
            data_re_out(0) => data_re_out(4),
            data_re_out(1) => data_re_out(36),
            data_re_out(2) => data_re_out(68),
            data_re_out(3) => data_re_out(100),
            data_re_out(4) => data_re_out(132),
            data_re_out(5) => data_re_out(164),
            data_re_out(6) => data_re_out(196),
            data_re_out(7) => data_re_out(228),
            data_re_out(8) => data_re_out(260),
            data_re_out(9) => data_re_out(292),
            data_re_out(10) => data_re_out(324),
            data_re_out(11) => data_re_out(356),
            data_re_out(12) => data_re_out(388),
            data_re_out(13) => data_re_out(420),
            data_re_out(14) => data_re_out(452),
            data_re_out(15) => data_re_out(484),
            data_re_out(16) => data_re_out(516),
            data_re_out(17) => data_re_out(548),
            data_re_out(18) => data_re_out(580),
            data_re_out(19) => data_re_out(612),
            data_re_out(20) => data_re_out(644),
            data_re_out(21) => data_re_out(676),
            data_re_out(22) => data_re_out(708),
            data_re_out(23) => data_re_out(740),
            data_re_out(24) => data_re_out(772),
            data_re_out(25) => data_re_out(804),
            data_re_out(26) => data_re_out(836),
            data_re_out(27) => data_re_out(868),
            data_re_out(28) => data_re_out(900),
            data_re_out(29) => data_re_out(932),
            data_re_out(30) => data_re_out(964),
            data_re_out(31) => data_re_out(996),
            data_re_out(32) => data_re_out(1028),
            data_re_out(33) => data_re_out(1060),
            data_re_out(34) => data_re_out(1092),
            data_re_out(35) => data_re_out(1124),
            data_re_out(36) => data_re_out(1156),
            data_re_out(37) => data_re_out(1188),
            data_re_out(38) => data_re_out(1220),
            data_re_out(39) => data_re_out(1252),
            data_re_out(40) => data_re_out(1284),
            data_re_out(41) => data_re_out(1316),
            data_re_out(42) => data_re_out(1348),
            data_re_out(43) => data_re_out(1380),
            data_re_out(44) => data_re_out(1412),
            data_re_out(45) => data_re_out(1444),
            data_re_out(46) => data_re_out(1476),
            data_re_out(47) => data_re_out(1508),
            data_re_out(48) => data_re_out(1540),
            data_re_out(49) => data_re_out(1572),
            data_re_out(50) => data_re_out(1604),
            data_re_out(51) => data_re_out(1636),
            data_re_out(52) => data_re_out(1668),
            data_re_out(53) => data_re_out(1700),
            data_re_out(54) => data_re_out(1732),
            data_re_out(55) => data_re_out(1764),
            data_re_out(56) => data_re_out(1796),
            data_re_out(57) => data_re_out(1828),
            data_re_out(58) => data_re_out(1860),
            data_re_out(59) => data_re_out(1892),
            data_re_out(60) => data_re_out(1924),
            data_re_out(61) => data_re_out(1956),
            data_re_out(62) => data_re_out(1988),
            data_re_out(63) => data_re_out(2020),
            data_im_out(0) => data_im_out(4),
            data_im_out(1) => data_im_out(36),
            data_im_out(2) => data_im_out(68),
            data_im_out(3) => data_im_out(100),
            data_im_out(4) => data_im_out(132),
            data_im_out(5) => data_im_out(164),
            data_im_out(6) => data_im_out(196),
            data_im_out(7) => data_im_out(228),
            data_im_out(8) => data_im_out(260),
            data_im_out(9) => data_im_out(292),
            data_im_out(10) => data_im_out(324),
            data_im_out(11) => data_im_out(356),
            data_im_out(12) => data_im_out(388),
            data_im_out(13) => data_im_out(420),
            data_im_out(14) => data_im_out(452),
            data_im_out(15) => data_im_out(484),
            data_im_out(16) => data_im_out(516),
            data_im_out(17) => data_im_out(548),
            data_im_out(18) => data_im_out(580),
            data_im_out(19) => data_im_out(612),
            data_im_out(20) => data_im_out(644),
            data_im_out(21) => data_im_out(676),
            data_im_out(22) => data_im_out(708),
            data_im_out(23) => data_im_out(740),
            data_im_out(24) => data_im_out(772),
            data_im_out(25) => data_im_out(804),
            data_im_out(26) => data_im_out(836),
            data_im_out(27) => data_im_out(868),
            data_im_out(28) => data_im_out(900),
            data_im_out(29) => data_im_out(932),
            data_im_out(30) => data_im_out(964),
            data_im_out(31) => data_im_out(996),
            data_im_out(32) => data_im_out(1028),
            data_im_out(33) => data_im_out(1060),
            data_im_out(34) => data_im_out(1092),
            data_im_out(35) => data_im_out(1124),
            data_im_out(36) => data_im_out(1156),
            data_im_out(37) => data_im_out(1188),
            data_im_out(38) => data_im_out(1220),
            data_im_out(39) => data_im_out(1252),
            data_im_out(40) => data_im_out(1284),
            data_im_out(41) => data_im_out(1316),
            data_im_out(42) => data_im_out(1348),
            data_im_out(43) => data_im_out(1380),
            data_im_out(44) => data_im_out(1412),
            data_im_out(45) => data_im_out(1444),
            data_im_out(46) => data_im_out(1476),
            data_im_out(47) => data_im_out(1508),
            data_im_out(48) => data_im_out(1540),
            data_im_out(49) => data_im_out(1572),
            data_im_out(50) => data_im_out(1604),
            data_im_out(51) => data_im_out(1636),
            data_im_out(52) => data_im_out(1668),
            data_im_out(53) => data_im_out(1700),
            data_im_out(54) => data_im_out(1732),
            data_im_out(55) => data_im_out(1764),
            data_im_out(56) => data_im_out(1796),
            data_im_out(57) => data_im_out(1828),
            data_im_out(58) => data_im_out(1860),
            data_im_out(59) => data_im_out(1892),
            data_im_out(60) => data_im_out(1924),
            data_im_out(61) => data_im_out(1956),
            data_im_out(62) => data_im_out(1988),
            data_im_out(63) => data_im_out(2020)
        );           

    URFFT_PT64_5 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(320),
            data_re_in(1) => mul_re_out(321),
            data_re_in(2) => mul_re_out(322),
            data_re_in(3) => mul_re_out(323),
            data_re_in(4) => mul_re_out(324),
            data_re_in(5) => mul_re_out(325),
            data_re_in(6) => mul_re_out(326),
            data_re_in(7) => mul_re_out(327),
            data_re_in(8) => mul_re_out(328),
            data_re_in(9) => mul_re_out(329),
            data_re_in(10) => mul_re_out(330),
            data_re_in(11) => mul_re_out(331),
            data_re_in(12) => mul_re_out(332),
            data_re_in(13) => mul_re_out(333),
            data_re_in(14) => mul_re_out(334),
            data_re_in(15) => mul_re_out(335),
            data_re_in(16) => mul_re_out(336),
            data_re_in(17) => mul_re_out(337),
            data_re_in(18) => mul_re_out(338),
            data_re_in(19) => mul_re_out(339),
            data_re_in(20) => mul_re_out(340),
            data_re_in(21) => mul_re_out(341),
            data_re_in(22) => mul_re_out(342),
            data_re_in(23) => mul_re_out(343),
            data_re_in(24) => mul_re_out(344),
            data_re_in(25) => mul_re_out(345),
            data_re_in(26) => mul_re_out(346),
            data_re_in(27) => mul_re_out(347),
            data_re_in(28) => mul_re_out(348),
            data_re_in(29) => mul_re_out(349),
            data_re_in(30) => mul_re_out(350),
            data_re_in(31) => mul_re_out(351),
            data_re_in(32) => mul_re_out(352),
            data_re_in(33) => mul_re_out(353),
            data_re_in(34) => mul_re_out(354),
            data_re_in(35) => mul_re_out(355),
            data_re_in(36) => mul_re_out(356),
            data_re_in(37) => mul_re_out(357),
            data_re_in(38) => mul_re_out(358),
            data_re_in(39) => mul_re_out(359),
            data_re_in(40) => mul_re_out(360),
            data_re_in(41) => mul_re_out(361),
            data_re_in(42) => mul_re_out(362),
            data_re_in(43) => mul_re_out(363),
            data_re_in(44) => mul_re_out(364),
            data_re_in(45) => mul_re_out(365),
            data_re_in(46) => mul_re_out(366),
            data_re_in(47) => mul_re_out(367),
            data_re_in(48) => mul_re_out(368),
            data_re_in(49) => mul_re_out(369),
            data_re_in(50) => mul_re_out(370),
            data_re_in(51) => mul_re_out(371),
            data_re_in(52) => mul_re_out(372),
            data_re_in(53) => mul_re_out(373),
            data_re_in(54) => mul_re_out(374),
            data_re_in(55) => mul_re_out(375),
            data_re_in(56) => mul_re_out(376),
            data_re_in(57) => mul_re_out(377),
            data_re_in(58) => mul_re_out(378),
            data_re_in(59) => mul_re_out(379),
            data_re_in(60) => mul_re_out(380),
            data_re_in(61) => mul_re_out(381),
            data_re_in(62) => mul_re_out(382),
            data_re_in(63) => mul_re_out(383),
            data_im_in(0) => mul_im_out(320),
            data_im_in(1) => mul_im_out(321),
            data_im_in(2) => mul_im_out(322),
            data_im_in(3) => mul_im_out(323),
            data_im_in(4) => mul_im_out(324),
            data_im_in(5) => mul_im_out(325),
            data_im_in(6) => mul_im_out(326),
            data_im_in(7) => mul_im_out(327),
            data_im_in(8) => mul_im_out(328),
            data_im_in(9) => mul_im_out(329),
            data_im_in(10) => mul_im_out(330),
            data_im_in(11) => mul_im_out(331),
            data_im_in(12) => mul_im_out(332),
            data_im_in(13) => mul_im_out(333),
            data_im_in(14) => mul_im_out(334),
            data_im_in(15) => mul_im_out(335),
            data_im_in(16) => mul_im_out(336),
            data_im_in(17) => mul_im_out(337),
            data_im_in(18) => mul_im_out(338),
            data_im_in(19) => mul_im_out(339),
            data_im_in(20) => mul_im_out(340),
            data_im_in(21) => mul_im_out(341),
            data_im_in(22) => mul_im_out(342),
            data_im_in(23) => mul_im_out(343),
            data_im_in(24) => mul_im_out(344),
            data_im_in(25) => mul_im_out(345),
            data_im_in(26) => mul_im_out(346),
            data_im_in(27) => mul_im_out(347),
            data_im_in(28) => mul_im_out(348),
            data_im_in(29) => mul_im_out(349),
            data_im_in(30) => mul_im_out(350),
            data_im_in(31) => mul_im_out(351),
            data_im_in(32) => mul_im_out(352),
            data_im_in(33) => mul_im_out(353),
            data_im_in(34) => mul_im_out(354),
            data_im_in(35) => mul_im_out(355),
            data_im_in(36) => mul_im_out(356),
            data_im_in(37) => mul_im_out(357),
            data_im_in(38) => mul_im_out(358),
            data_im_in(39) => mul_im_out(359),
            data_im_in(40) => mul_im_out(360),
            data_im_in(41) => mul_im_out(361),
            data_im_in(42) => mul_im_out(362),
            data_im_in(43) => mul_im_out(363),
            data_im_in(44) => mul_im_out(364),
            data_im_in(45) => mul_im_out(365),
            data_im_in(46) => mul_im_out(366),
            data_im_in(47) => mul_im_out(367),
            data_im_in(48) => mul_im_out(368),
            data_im_in(49) => mul_im_out(369),
            data_im_in(50) => mul_im_out(370),
            data_im_in(51) => mul_im_out(371),
            data_im_in(52) => mul_im_out(372),
            data_im_in(53) => mul_im_out(373),
            data_im_in(54) => mul_im_out(374),
            data_im_in(55) => mul_im_out(375),
            data_im_in(56) => mul_im_out(376),
            data_im_in(57) => mul_im_out(377),
            data_im_in(58) => mul_im_out(378),
            data_im_in(59) => mul_im_out(379),
            data_im_in(60) => mul_im_out(380),
            data_im_in(61) => mul_im_out(381),
            data_im_in(62) => mul_im_out(382),
            data_im_in(63) => mul_im_out(383),
            data_re_out(0) => data_re_out(5),
            data_re_out(1) => data_re_out(37),
            data_re_out(2) => data_re_out(69),
            data_re_out(3) => data_re_out(101),
            data_re_out(4) => data_re_out(133),
            data_re_out(5) => data_re_out(165),
            data_re_out(6) => data_re_out(197),
            data_re_out(7) => data_re_out(229),
            data_re_out(8) => data_re_out(261),
            data_re_out(9) => data_re_out(293),
            data_re_out(10) => data_re_out(325),
            data_re_out(11) => data_re_out(357),
            data_re_out(12) => data_re_out(389),
            data_re_out(13) => data_re_out(421),
            data_re_out(14) => data_re_out(453),
            data_re_out(15) => data_re_out(485),
            data_re_out(16) => data_re_out(517),
            data_re_out(17) => data_re_out(549),
            data_re_out(18) => data_re_out(581),
            data_re_out(19) => data_re_out(613),
            data_re_out(20) => data_re_out(645),
            data_re_out(21) => data_re_out(677),
            data_re_out(22) => data_re_out(709),
            data_re_out(23) => data_re_out(741),
            data_re_out(24) => data_re_out(773),
            data_re_out(25) => data_re_out(805),
            data_re_out(26) => data_re_out(837),
            data_re_out(27) => data_re_out(869),
            data_re_out(28) => data_re_out(901),
            data_re_out(29) => data_re_out(933),
            data_re_out(30) => data_re_out(965),
            data_re_out(31) => data_re_out(997),
            data_re_out(32) => data_re_out(1029),
            data_re_out(33) => data_re_out(1061),
            data_re_out(34) => data_re_out(1093),
            data_re_out(35) => data_re_out(1125),
            data_re_out(36) => data_re_out(1157),
            data_re_out(37) => data_re_out(1189),
            data_re_out(38) => data_re_out(1221),
            data_re_out(39) => data_re_out(1253),
            data_re_out(40) => data_re_out(1285),
            data_re_out(41) => data_re_out(1317),
            data_re_out(42) => data_re_out(1349),
            data_re_out(43) => data_re_out(1381),
            data_re_out(44) => data_re_out(1413),
            data_re_out(45) => data_re_out(1445),
            data_re_out(46) => data_re_out(1477),
            data_re_out(47) => data_re_out(1509),
            data_re_out(48) => data_re_out(1541),
            data_re_out(49) => data_re_out(1573),
            data_re_out(50) => data_re_out(1605),
            data_re_out(51) => data_re_out(1637),
            data_re_out(52) => data_re_out(1669),
            data_re_out(53) => data_re_out(1701),
            data_re_out(54) => data_re_out(1733),
            data_re_out(55) => data_re_out(1765),
            data_re_out(56) => data_re_out(1797),
            data_re_out(57) => data_re_out(1829),
            data_re_out(58) => data_re_out(1861),
            data_re_out(59) => data_re_out(1893),
            data_re_out(60) => data_re_out(1925),
            data_re_out(61) => data_re_out(1957),
            data_re_out(62) => data_re_out(1989),
            data_re_out(63) => data_re_out(2021),
            data_im_out(0) => data_im_out(5),
            data_im_out(1) => data_im_out(37),
            data_im_out(2) => data_im_out(69),
            data_im_out(3) => data_im_out(101),
            data_im_out(4) => data_im_out(133),
            data_im_out(5) => data_im_out(165),
            data_im_out(6) => data_im_out(197),
            data_im_out(7) => data_im_out(229),
            data_im_out(8) => data_im_out(261),
            data_im_out(9) => data_im_out(293),
            data_im_out(10) => data_im_out(325),
            data_im_out(11) => data_im_out(357),
            data_im_out(12) => data_im_out(389),
            data_im_out(13) => data_im_out(421),
            data_im_out(14) => data_im_out(453),
            data_im_out(15) => data_im_out(485),
            data_im_out(16) => data_im_out(517),
            data_im_out(17) => data_im_out(549),
            data_im_out(18) => data_im_out(581),
            data_im_out(19) => data_im_out(613),
            data_im_out(20) => data_im_out(645),
            data_im_out(21) => data_im_out(677),
            data_im_out(22) => data_im_out(709),
            data_im_out(23) => data_im_out(741),
            data_im_out(24) => data_im_out(773),
            data_im_out(25) => data_im_out(805),
            data_im_out(26) => data_im_out(837),
            data_im_out(27) => data_im_out(869),
            data_im_out(28) => data_im_out(901),
            data_im_out(29) => data_im_out(933),
            data_im_out(30) => data_im_out(965),
            data_im_out(31) => data_im_out(997),
            data_im_out(32) => data_im_out(1029),
            data_im_out(33) => data_im_out(1061),
            data_im_out(34) => data_im_out(1093),
            data_im_out(35) => data_im_out(1125),
            data_im_out(36) => data_im_out(1157),
            data_im_out(37) => data_im_out(1189),
            data_im_out(38) => data_im_out(1221),
            data_im_out(39) => data_im_out(1253),
            data_im_out(40) => data_im_out(1285),
            data_im_out(41) => data_im_out(1317),
            data_im_out(42) => data_im_out(1349),
            data_im_out(43) => data_im_out(1381),
            data_im_out(44) => data_im_out(1413),
            data_im_out(45) => data_im_out(1445),
            data_im_out(46) => data_im_out(1477),
            data_im_out(47) => data_im_out(1509),
            data_im_out(48) => data_im_out(1541),
            data_im_out(49) => data_im_out(1573),
            data_im_out(50) => data_im_out(1605),
            data_im_out(51) => data_im_out(1637),
            data_im_out(52) => data_im_out(1669),
            data_im_out(53) => data_im_out(1701),
            data_im_out(54) => data_im_out(1733),
            data_im_out(55) => data_im_out(1765),
            data_im_out(56) => data_im_out(1797),
            data_im_out(57) => data_im_out(1829),
            data_im_out(58) => data_im_out(1861),
            data_im_out(59) => data_im_out(1893),
            data_im_out(60) => data_im_out(1925),
            data_im_out(61) => data_im_out(1957),
            data_im_out(62) => data_im_out(1989),
            data_im_out(63) => data_im_out(2021)
        );           

    URFFT_PT64_6 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(384),
            data_re_in(1) => mul_re_out(385),
            data_re_in(2) => mul_re_out(386),
            data_re_in(3) => mul_re_out(387),
            data_re_in(4) => mul_re_out(388),
            data_re_in(5) => mul_re_out(389),
            data_re_in(6) => mul_re_out(390),
            data_re_in(7) => mul_re_out(391),
            data_re_in(8) => mul_re_out(392),
            data_re_in(9) => mul_re_out(393),
            data_re_in(10) => mul_re_out(394),
            data_re_in(11) => mul_re_out(395),
            data_re_in(12) => mul_re_out(396),
            data_re_in(13) => mul_re_out(397),
            data_re_in(14) => mul_re_out(398),
            data_re_in(15) => mul_re_out(399),
            data_re_in(16) => mul_re_out(400),
            data_re_in(17) => mul_re_out(401),
            data_re_in(18) => mul_re_out(402),
            data_re_in(19) => mul_re_out(403),
            data_re_in(20) => mul_re_out(404),
            data_re_in(21) => mul_re_out(405),
            data_re_in(22) => mul_re_out(406),
            data_re_in(23) => mul_re_out(407),
            data_re_in(24) => mul_re_out(408),
            data_re_in(25) => mul_re_out(409),
            data_re_in(26) => mul_re_out(410),
            data_re_in(27) => mul_re_out(411),
            data_re_in(28) => mul_re_out(412),
            data_re_in(29) => mul_re_out(413),
            data_re_in(30) => mul_re_out(414),
            data_re_in(31) => mul_re_out(415),
            data_re_in(32) => mul_re_out(416),
            data_re_in(33) => mul_re_out(417),
            data_re_in(34) => mul_re_out(418),
            data_re_in(35) => mul_re_out(419),
            data_re_in(36) => mul_re_out(420),
            data_re_in(37) => mul_re_out(421),
            data_re_in(38) => mul_re_out(422),
            data_re_in(39) => mul_re_out(423),
            data_re_in(40) => mul_re_out(424),
            data_re_in(41) => mul_re_out(425),
            data_re_in(42) => mul_re_out(426),
            data_re_in(43) => mul_re_out(427),
            data_re_in(44) => mul_re_out(428),
            data_re_in(45) => mul_re_out(429),
            data_re_in(46) => mul_re_out(430),
            data_re_in(47) => mul_re_out(431),
            data_re_in(48) => mul_re_out(432),
            data_re_in(49) => mul_re_out(433),
            data_re_in(50) => mul_re_out(434),
            data_re_in(51) => mul_re_out(435),
            data_re_in(52) => mul_re_out(436),
            data_re_in(53) => mul_re_out(437),
            data_re_in(54) => mul_re_out(438),
            data_re_in(55) => mul_re_out(439),
            data_re_in(56) => mul_re_out(440),
            data_re_in(57) => mul_re_out(441),
            data_re_in(58) => mul_re_out(442),
            data_re_in(59) => mul_re_out(443),
            data_re_in(60) => mul_re_out(444),
            data_re_in(61) => mul_re_out(445),
            data_re_in(62) => mul_re_out(446),
            data_re_in(63) => mul_re_out(447),
            data_im_in(0) => mul_im_out(384),
            data_im_in(1) => mul_im_out(385),
            data_im_in(2) => mul_im_out(386),
            data_im_in(3) => mul_im_out(387),
            data_im_in(4) => mul_im_out(388),
            data_im_in(5) => mul_im_out(389),
            data_im_in(6) => mul_im_out(390),
            data_im_in(7) => mul_im_out(391),
            data_im_in(8) => mul_im_out(392),
            data_im_in(9) => mul_im_out(393),
            data_im_in(10) => mul_im_out(394),
            data_im_in(11) => mul_im_out(395),
            data_im_in(12) => mul_im_out(396),
            data_im_in(13) => mul_im_out(397),
            data_im_in(14) => mul_im_out(398),
            data_im_in(15) => mul_im_out(399),
            data_im_in(16) => mul_im_out(400),
            data_im_in(17) => mul_im_out(401),
            data_im_in(18) => mul_im_out(402),
            data_im_in(19) => mul_im_out(403),
            data_im_in(20) => mul_im_out(404),
            data_im_in(21) => mul_im_out(405),
            data_im_in(22) => mul_im_out(406),
            data_im_in(23) => mul_im_out(407),
            data_im_in(24) => mul_im_out(408),
            data_im_in(25) => mul_im_out(409),
            data_im_in(26) => mul_im_out(410),
            data_im_in(27) => mul_im_out(411),
            data_im_in(28) => mul_im_out(412),
            data_im_in(29) => mul_im_out(413),
            data_im_in(30) => mul_im_out(414),
            data_im_in(31) => mul_im_out(415),
            data_im_in(32) => mul_im_out(416),
            data_im_in(33) => mul_im_out(417),
            data_im_in(34) => mul_im_out(418),
            data_im_in(35) => mul_im_out(419),
            data_im_in(36) => mul_im_out(420),
            data_im_in(37) => mul_im_out(421),
            data_im_in(38) => mul_im_out(422),
            data_im_in(39) => mul_im_out(423),
            data_im_in(40) => mul_im_out(424),
            data_im_in(41) => mul_im_out(425),
            data_im_in(42) => mul_im_out(426),
            data_im_in(43) => mul_im_out(427),
            data_im_in(44) => mul_im_out(428),
            data_im_in(45) => mul_im_out(429),
            data_im_in(46) => mul_im_out(430),
            data_im_in(47) => mul_im_out(431),
            data_im_in(48) => mul_im_out(432),
            data_im_in(49) => mul_im_out(433),
            data_im_in(50) => mul_im_out(434),
            data_im_in(51) => mul_im_out(435),
            data_im_in(52) => mul_im_out(436),
            data_im_in(53) => mul_im_out(437),
            data_im_in(54) => mul_im_out(438),
            data_im_in(55) => mul_im_out(439),
            data_im_in(56) => mul_im_out(440),
            data_im_in(57) => mul_im_out(441),
            data_im_in(58) => mul_im_out(442),
            data_im_in(59) => mul_im_out(443),
            data_im_in(60) => mul_im_out(444),
            data_im_in(61) => mul_im_out(445),
            data_im_in(62) => mul_im_out(446),
            data_im_in(63) => mul_im_out(447),
            data_re_out(0) => data_re_out(6),
            data_re_out(1) => data_re_out(38),
            data_re_out(2) => data_re_out(70),
            data_re_out(3) => data_re_out(102),
            data_re_out(4) => data_re_out(134),
            data_re_out(5) => data_re_out(166),
            data_re_out(6) => data_re_out(198),
            data_re_out(7) => data_re_out(230),
            data_re_out(8) => data_re_out(262),
            data_re_out(9) => data_re_out(294),
            data_re_out(10) => data_re_out(326),
            data_re_out(11) => data_re_out(358),
            data_re_out(12) => data_re_out(390),
            data_re_out(13) => data_re_out(422),
            data_re_out(14) => data_re_out(454),
            data_re_out(15) => data_re_out(486),
            data_re_out(16) => data_re_out(518),
            data_re_out(17) => data_re_out(550),
            data_re_out(18) => data_re_out(582),
            data_re_out(19) => data_re_out(614),
            data_re_out(20) => data_re_out(646),
            data_re_out(21) => data_re_out(678),
            data_re_out(22) => data_re_out(710),
            data_re_out(23) => data_re_out(742),
            data_re_out(24) => data_re_out(774),
            data_re_out(25) => data_re_out(806),
            data_re_out(26) => data_re_out(838),
            data_re_out(27) => data_re_out(870),
            data_re_out(28) => data_re_out(902),
            data_re_out(29) => data_re_out(934),
            data_re_out(30) => data_re_out(966),
            data_re_out(31) => data_re_out(998),
            data_re_out(32) => data_re_out(1030),
            data_re_out(33) => data_re_out(1062),
            data_re_out(34) => data_re_out(1094),
            data_re_out(35) => data_re_out(1126),
            data_re_out(36) => data_re_out(1158),
            data_re_out(37) => data_re_out(1190),
            data_re_out(38) => data_re_out(1222),
            data_re_out(39) => data_re_out(1254),
            data_re_out(40) => data_re_out(1286),
            data_re_out(41) => data_re_out(1318),
            data_re_out(42) => data_re_out(1350),
            data_re_out(43) => data_re_out(1382),
            data_re_out(44) => data_re_out(1414),
            data_re_out(45) => data_re_out(1446),
            data_re_out(46) => data_re_out(1478),
            data_re_out(47) => data_re_out(1510),
            data_re_out(48) => data_re_out(1542),
            data_re_out(49) => data_re_out(1574),
            data_re_out(50) => data_re_out(1606),
            data_re_out(51) => data_re_out(1638),
            data_re_out(52) => data_re_out(1670),
            data_re_out(53) => data_re_out(1702),
            data_re_out(54) => data_re_out(1734),
            data_re_out(55) => data_re_out(1766),
            data_re_out(56) => data_re_out(1798),
            data_re_out(57) => data_re_out(1830),
            data_re_out(58) => data_re_out(1862),
            data_re_out(59) => data_re_out(1894),
            data_re_out(60) => data_re_out(1926),
            data_re_out(61) => data_re_out(1958),
            data_re_out(62) => data_re_out(1990),
            data_re_out(63) => data_re_out(2022),
            data_im_out(0) => data_im_out(6),
            data_im_out(1) => data_im_out(38),
            data_im_out(2) => data_im_out(70),
            data_im_out(3) => data_im_out(102),
            data_im_out(4) => data_im_out(134),
            data_im_out(5) => data_im_out(166),
            data_im_out(6) => data_im_out(198),
            data_im_out(7) => data_im_out(230),
            data_im_out(8) => data_im_out(262),
            data_im_out(9) => data_im_out(294),
            data_im_out(10) => data_im_out(326),
            data_im_out(11) => data_im_out(358),
            data_im_out(12) => data_im_out(390),
            data_im_out(13) => data_im_out(422),
            data_im_out(14) => data_im_out(454),
            data_im_out(15) => data_im_out(486),
            data_im_out(16) => data_im_out(518),
            data_im_out(17) => data_im_out(550),
            data_im_out(18) => data_im_out(582),
            data_im_out(19) => data_im_out(614),
            data_im_out(20) => data_im_out(646),
            data_im_out(21) => data_im_out(678),
            data_im_out(22) => data_im_out(710),
            data_im_out(23) => data_im_out(742),
            data_im_out(24) => data_im_out(774),
            data_im_out(25) => data_im_out(806),
            data_im_out(26) => data_im_out(838),
            data_im_out(27) => data_im_out(870),
            data_im_out(28) => data_im_out(902),
            data_im_out(29) => data_im_out(934),
            data_im_out(30) => data_im_out(966),
            data_im_out(31) => data_im_out(998),
            data_im_out(32) => data_im_out(1030),
            data_im_out(33) => data_im_out(1062),
            data_im_out(34) => data_im_out(1094),
            data_im_out(35) => data_im_out(1126),
            data_im_out(36) => data_im_out(1158),
            data_im_out(37) => data_im_out(1190),
            data_im_out(38) => data_im_out(1222),
            data_im_out(39) => data_im_out(1254),
            data_im_out(40) => data_im_out(1286),
            data_im_out(41) => data_im_out(1318),
            data_im_out(42) => data_im_out(1350),
            data_im_out(43) => data_im_out(1382),
            data_im_out(44) => data_im_out(1414),
            data_im_out(45) => data_im_out(1446),
            data_im_out(46) => data_im_out(1478),
            data_im_out(47) => data_im_out(1510),
            data_im_out(48) => data_im_out(1542),
            data_im_out(49) => data_im_out(1574),
            data_im_out(50) => data_im_out(1606),
            data_im_out(51) => data_im_out(1638),
            data_im_out(52) => data_im_out(1670),
            data_im_out(53) => data_im_out(1702),
            data_im_out(54) => data_im_out(1734),
            data_im_out(55) => data_im_out(1766),
            data_im_out(56) => data_im_out(1798),
            data_im_out(57) => data_im_out(1830),
            data_im_out(58) => data_im_out(1862),
            data_im_out(59) => data_im_out(1894),
            data_im_out(60) => data_im_out(1926),
            data_im_out(61) => data_im_out(1958),
            data_im_out(62) => data_im_out(1990),
            data_im_out(63) => data_im_out(2022)
        );           

    URFFT_PT64_7 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(448),
            data_re_in(1) => mul_re_out(449),
            data_re_in(2) => mul_re_out(450),
            data_re_in(3) => mul_re_out(451),
            data_re_in(4) => mul_re_out(452),
            data_re_in(5) => mul_re_out(453),
            data_re_in(6) => mul_re_out(454),
            data_re_in(7) => mul_re_out(455),
            data_re_in(8) => mul_re_out(456),
            data_re_in(9) => mul_re_out(457),
            data_re_in(10) => mul_re_out(458),
            data_re_in(11) => mul_re_out(459),
            data_re_in(12) => mul_re_out(460),
            data_re_in(13) => mul_re_out(461),
            data_re_in(14) => mul_re_out(462),
            data_re_in(15) => mul_re_out(463),
            data_re_in(16) => mul_re_out(464),
            data_re_in(17) => mul_re_out(465),
            data_re_in(18) => mul_re_out(466),
            data_re_in(19) => mul_re_out(467),
            data_re_in(20) => mul_re_out(468),
            data_re_in(21) => mul_re_out(469),
            data_re_in(22) => mul_re_out(470),
            data_re_in(23) => mul_re_out(471),
            data_re_in(24) => mul_re_out(472),
            data_re_in(25) => mul_re_out(473),
            data_re_in(26) => mul_re_out(474),
            data_re_in(27) => mul_re_out(475),
            data_re_in(28) => mul_re_out(476),
            data_re_in(29) => mul_re_out(477),
            data_re_in(30) => mul_re_out(478),
            data_re_in(31) => mul_re_out(479),
            data_re_in(32) => mul_re_out(480),
            data_re_in(33) => mul_re_out(481),
            data_re_in(34) => mul_re_out(482),
            data_re_in(35) => mul_re_out(483),
            data_re_in(36) => mul_re_out(484),
            data_re_in(37) => mul_re_out(485),
            data_re_in(38) => mul_re_out(486),
            data_re_in(39) => mul_re_out(487),
            data_re_in(40) => mul_re_out(488),
            data_re_in(41) => mul_re_out(489),
            data_re_in(42) => mul_re_out(490),
            data_re_in(43) => mul_re_out(491),
            data_re_in(44) => mul_re_out(492),
            data_re_in(45) => mul_re_out(493),
            data_re_in(46) => mul_re_out(494),
            data_re_in(47) => mul_re_out(495),
            data_re_in(48) => mul_re_out(496),
            data_re_in(49) => mul_re_out(497),
            data_re_in(50) => mul_re_out(498),
            data_re_in(51) => mul_re_out(499),
            data_re_in(52) => mul_re_out(500),
            data_re_in(53) => mul_re_out(501),
            data_re_in(54) => mul_re_out(502),
            data_re_in(55) => mul_re_out(503),
            data_re_in(56) => mul_re_out(504),
            data_re_in(57) => mul_re_out(505),
            data_re_in(58) => mul_re_out(506),
            data_re_in(59) => mul_re_out(507),
            data_re_in(60) => mul_re_out(508),
            data_re_in(61) => mul_re_out(509),
            data_re_in(62) => mul_re_out(510),
            data_re_in(63) => mul_re_out(511),
            data_im_in(0) => mul_im_out(448),
            data_im_in(1) => mul_im_out(449),
            data_im_in(2) => mul_im_out(450),
            data_im_in(3) => mul_im_out(451),
            data_im_in(4) => mul_im_out(452),
            data_im_in(5) => mul_im_out(453),
            data_im_in(6) => mul_im_out(454),
            data_im_in(7) => mul_im_out(455),
            data_im_in(8) => mul_im_out(456),
            data_im_in(9) => mul_im_out(457),
            data_im_in(10) => mul_im_out(458),
            data_im_in(11) => mul_im_out(459),
            data_im_in(12) => mul_im_out(460),
            data_im_in(13) => mul_im_out(461),
            data_im_in(14) => mul_im_out(462),
            data_im_in(15) => mul_im_out(463),
            data_im_in(16) => mul_im_out(464),
            data_im_in(17) => mul_im_out(465),
            data_im_in(18) => mul_im_out(466),
            data_im_in(19) => mul_im_out(467),
            data_im_in(20) => mul_im_out(468),
            data_im_in(21) => mul_im_out(469),
            data_im_in(22) => mul_im_out(470),
            data_im_in(23) => mul_im_out(471),
            data_im_in(24) => mul_im_out(472),
            data_im_in(25) => mul_im_out(473),
            data_im_in(26) => mul_im_out(474),
            data_im_in(27) => mul_im_out(475),
            data_im_in(28) => mul_im_out(476),
            data_im_in(29) => mul_im_out(477),
            data_im_in(30) => mul_im_out(478),
            data_im_in(31) => mul_im_out(479),
            data_im_in(32) => mul_im_out(480),
            data_im_in(33) => mul_im_out(481),
            data_im_in(34) => mul_im_out(482),
            data_im_in(35) => mul_im_out(483),
            data_im_in(36) => mul_im_out(484),
            data_im_in(37) => mul_im_out(485),
            data_im_in(38) => mul_im_out(486),
            data_im_in(39) => mul_im_out(487),
            data_im_in(40) => mul_im_out(488),
            data_im_in(41) => mul_im_out(489),
            data_im_in(42) => mul_im_out(490),
            data_im_in(43) => mul_im_out(491),
            data_im_in(44) => mul_im_out(492),
            data_im_in(45) => mul_im_out(493),
            data_im_in(46) => mul_im_out(494),
            data_im_in(47) => mul_im_out(495),
            data_im_in(48) => mul_im_out(496),
            data_im_in(49) => mul_im_out(497),
            data_im_in(50) => mul_im_out(498),
            data_im_in(51) => mul_im_out(499),
            data_im_in(52) => mul_im_out(500),
            data_im_in(53) => mul_im_out(501),
            data_im_in(54) => mul_im_out(502),
            data_im_in(55) => mul_im_out(503),
            data_im_in(56) => mul_im_out(504),
            data_im_in(57) => mul_im_out(505),
            data_im_in(58) => mul_im_out(506),
            data_im_in(59) => mul_im_out(507),
            data_im_in(60) => mul_im_out(508),
            data_im_in(61) => mul_im_out(509),
            data_im_in(62) => mul_im_out(510),
            data_im_in(63) => mul_im_out(511),
            data_re_out(0) => data_re_out(7),
            data_re_out(1) => data_re_out(39),
            data_re_out(2) => data_re_out(71),
            data_re_out(3) => data_re_out(103),
            data_re_out(4) => data_re_out(135),
            data_re_out(5) => data_re_out(167),
            data_re_out(6) => data_re_out(199),
            data_re_out(7) => data_re_out(231),
            data_re_out(8) => data_re_out(263),
            data_re_out(9) => data_re_out(295),
            data_re_out(10) => data_re_out(327),
            data_re_out(11) => data_re_out(359),
            data_re_out(12) => data_re_out(391),
            data_re_out(13) => data_re_out(423),
            data_re_out(14) => data_re_out(455),
            data_re_out(15) => data_re_out(487),
            data_re_out(16) => data_re_out(519),
            data_re_out(17) => data_re_out(551),
            data_re_out(18) => data_re_out(583),
            data_re_out(19) => data_re_out(615),
            data_re_out(20) => data_re_out(647),
            data_re_out(21) => data_re_out(679),
            data_re_out(22) => data_re_out(711),
            data_re_out(23) => data_re_out(743),
            data_re_out(24) => data_re_out(775),
            data_re_out(25) => data_re_out(807),
            data_re_out(26) => data_re_out(839),
            data_re_out(27) => data_re_out(871),
            data_re_out(28) => data_re_out(903),
            data_re_out(29) => data_re_out(935),
            data_re_out(30) => data_re_out(967),
            data_re_out(31) => data_re_out(999),
            data_re_out(32) => data_re_out(1031),
            data_re_out(33) => data_re_out(1063),
            data_re_out(34) => data_re_out(1095),
            data_re_out(35) => data_re_out(1127),
            data_re_out(36) => data_re_out(1159),
            data_re_out(37) => data_re_out(1191),
            data_re_out(38) => data_re_out(1223),
            data_re_out(39) => data_re_out(1255),
            data_re_out(40) => data_re_out(1287),
            data_re_out(41) => data_re_out(1319),
            data_re_out(42) => data_re_out(1351),
            data_re_out(43) => data_re_out(1383),
            data_re_out(44) => data_re_out(1415),
            data_re_out(45) => data_re_out(1447),
            data_re_out(46) => data_re_out(1479),
            data_re_out(47) => data_re_out(1511),
            data_re_out(48) => data_re_out(1543),
            data_re_out(49) => data_re_out(1575),
            data_re_out(50) => data_re_out(1607),
            data_re_out(51) => data_re_out(1639),
            data_re_out(52) => data_re_out(1671),
            data_re_out(53) => data_re_out(1703),
            data_re_out(54) => data_re_out(1735),
            data_re_out(55) => data_re_out(1767),
            data_re_out(56) => data_re_out(1799),
            data_re_out(57) => data_re_out(1831),
            data_re_out(58) => data_re_out(1863),
            data_re_out(59) => data_re_out(1895),
            data_re_out(60) => data_re_out(1927),
            data_re_out(61) => data_re_out(1959),
            data_re_out(62) => data_re_out(1991),
            data_re_out(63) => data_re_out(2023),
            data_im_out(0) => data_im_out(7),
            data_im_out(1) => data_im_out(39),
            data_im_out(2) => data_im_out(71),
            data_im_out(3) => data_im_out(103),
            data_im_out(4) => data_im_out(135),
            data_im_out(5) => data_im_out(167),
            data_im_out(6) => data_im_out(199),
            data_im_out(7) => data_im_out(231),
            data_im_out(8) => data_im_out(263),
            data_im_out(9) => data_im_out(295),
            data_im_out(10) => data_im_out(327),
            data_im_out(11) => data_im_out(359),
            data_im_out(12) => data_im_out(391),
            data_im_out(13) => data_im_out(423),
            data_im_out(14) => data_im_out(455),
            data_im_out(15) => data_im_out(487),
            data_im_out(16) => data_im_out(519),
            data_im_out(17) => data_im_out(551),
            data_im_out(18) => data_im_out(583),
            data_im_out(19) => data_im_out(615),
            data_im_out(20) => data_im_out(647),
            data_im_out(21) => data_im_out(679),
            data_im_out(22) => data_im_out(711),
            data_im_out(23) => data_im_out(743),
            data_im_out(24) => data_im_out(775),
            data_im_out(25) => data_im_out(807),
            data_im_out(26) => data_im_out(839),
            data_im_out(27) => data_im_out(871),
            data_im_out(28) => data_im_out(903),
            data_im_out(29) => data_im_out(935),
            data_im_out(30) => data_im_out(967),
            data_im_out(31) => data_im_out(999),
            data_im_out(32) => data_im_out(1031),
            data_im_out(33) => data_im_out(1063),
            data_im_out(34) => data_im_out(1095),
            data_im_out(35) => data_im_out(1127),
            data_im_out(36) => data_im_out(1159),
            data_im_out(37) => data_im_out(1191),
            data_im_out(38) => data_im_out(1223),
            data_im_out(39) => data_im_out(1255),
            data_im_out(40) => data_im_out(1287),
            data_im_out(41) => data_im_out(1319),
            data_im_out(42) => data_im_out(1351),
            data_im_out(43) => data_im_out(1383),
            data_im_out(44) => data_im_out(1415),
            data_im_out(45) => data_im_out(1447),
            data_im_out(46) => data_im_out(1479),
            data_im_out(47) => data_im_out(1511),
            data_im_out(48) => data_im_out(1543),
            data_im_out(49) => data_im_out(1575),
            data_im_out(50) => data_im_out(1607),
            data_im_out(51) => data_im_out(1639),
            data_im_out(52) => data_im_out(1671),
            data_im_out(53) => data_im_out(1703),
            data_im_out(54) => data_im_out(1735),
            data_im_out(55) => data_im_out(1767),
            data_im_out(56) => data_im_out(1799),
            data_im_out(57) => data_im_out(1831),
            data_im_out(58) => data_im_out(1863),
            data_im_out(59) => data_im_out(1895),
            data_im_out(60) => data_im_out(1927),
            data_im_out(61) => data_im_out(1959),
            data_im_out(62) => data_im_out(1991),
            data_im_out(63) => data_im_out(2023)
        );           

    URFFT_PT64_8 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(512),
            data_re_in(1) => mul_re_out(513),
            data_re_in(2) => mul_re_out(514),
            data_re_in(3) => mul_re_out(515),
            data_re_in(4) => mul_re_out(516),
            data_re_in(5) => mul_re_out(517),
            data_re_in(6) => mul_re_out(518),
            data_re_in(7) => mul_re_out(519),
            data_re_in(8) => mul_re_out(520),
            data_re_in(9) => mul_re_out(521),
            data_re_in(10) => mul_re_out(522),
            data_re_in(11) => mul_re_out(523),
            data_re_in(12) => mul_re_out(524),
            data_re_in(13) => mul_re_out(525),
            data_re_in(14) => mul_re_out(526),
            data_re_in(15) => mul_re_out(527),
            data_re_in(16) => mul_re_out(528),
            data_re_in(17) => mul_re_out(529),
            data_re_in(18) => mul_re_out(530),
            data_re_in(19) => mul_re_out(531),
            data_re_in(20) => mul_re_out(532),
            data_re_in(21) => mul_re_out(533),
            data_re_in(22) => mul_re_out(534),
            data_re_in(23) => mul_re_out(535),
            data_re_in(24) => mul_re_out(536),
            data_re_in(25) => mul_re_out(537),
            data_re_in(26) => mul_re_out(538),
            data_re_in(27) => mul_re_out(539),
            data_re_in(28) => mul_re_out(540),
            data_re_in(29) => mul_re_out(541),
            data_re_in(30) => mul_re_out(542),
            data_re_in(31) => mul_re_out(543),
            data_re_in(32) => mul_re_out(544),
            data_re_in(33) => mul_re_out(545),
            data_re_in(34) => mul_re_out(546),
            data_re_in(35) => mul_re_out(547),
            data_re_in(36) => mul_re_out(548),
            data_re_in(37) => mul_re_out(549),
            data_re_in(38) => mul_re_out(550),
            data_re_in(39) => mul_re_out(551),
            data_re_in(40) => mul_re_out(552),
            data_re_in(41) => mul_re_out(553),
            data_re_in(42) => mul_re_out(554),
            data_re_in(43) => mul_re_out(555),
            data_re_in(44) => mul_re_out(556),
            data_re_in(45) => mul_re_out(557),
            data_re_in(46) => mul_re_out(558),
            data_re_in(47) => mul_re_out(559),
            data_re_in(48) => mul_re_out(560),
            data_re_in(49) => mul_re_out(561),
            data_re_in(50) => mul_re_out(562),
            data_re_in(51) => mul_re_out(563),
            data_re_in(52) => mul_re_out(564),
            data_re_in(53) => mul_re_out(565),
            data_re_in(54) => mul_re_out(566),
            data_re_in(55) => mul_re_out(567),
            data_re_in(56) => mul_re_out(568),
            data_re_in(57) => mul_re_out(569),
            data_re_in(58) => mul_re_out(570),
            data_re_in(59) => mul_re_out(571),
            data_re_in(60) => mul_re_out(572),
            data_re_in(61) => mul_re_out(573),
            data_re_in(62) => mul_re_out(574),
            data_re_in(63) => mul_re_out(575),
            data_im_in(0) => mul_im_out(512),
            data_im_in(1) => mul_im_out(513),
            data_im_in(2) => mul_im_out(514),
            data_im_in(3) => mul_im_out(515),
            data_im_in(4) => mul_im_out(516),
            data_im_in(5) => mul_im_out(517),
            data_im_in(6) => mul_im_out(518),
            data_im_in(7) => mul_im_out(519),
            data_im_in(8) => mul_im_out(520),
            data_im_in(9) => mul_im_out(521),
            data_im_in(10) => mul_im_out(522),
            data_im_in(11) => mul_im_out(523),
            data_im_in(12) => mul_im_out(524),
            data_im_in(13) => mul_im_out(525),
            data_im_in(14) => mul_im_out(526),
            data_im_in(15) => mul_im_out(527),
            data_im_in(16) => mul_im_out(528),
            data_im_in(17) => mul_im_out(529),
            data_im_in(18) => mul_im_out(530),
            data_im_in(19) => mul_im_out(531),
            data_im_in(20) => mul_im_out(532),
            data_im_in(21) => mul_im_out(533),
            data_im_in(22) => mul_im_out(534),
            data_im_in(23) => mul_im_out(535),
            data_im_in(24) => mul_im_out(536),
            data_im_in(25) => mul_im_out(537),
            data_im_in(26) => mul_im_out(538),
            data_im_in(27) => mul_im_out(539),
            data_im_in(28) => mul_im_out(540),
            data_im_in(29) => mul_im_out(541),
            data_im_in(30) => mul_im_out(542),
            data_im_in(31) => mul_im_out(543),
            data_im_in(32) => mul_im_out(544),
            data_im_in(33) => mul_im_out(545),
            data_im_in(34) => mul_im_out(546),
            data_im_in(35) => mul_im_out(547),
            data_im_in(36) => mul_im_out(548),
            data_im_in(37) => mul_im_out(549),
            data_im_in(38) => mul_im_out(550),
            data_im_in(39) => mul_im_out(551),
            data_im_in(40) => mul_im_out(552),
            data_im_in(41) => mul_im_out(553),
            data_im_in(42) => mul_im_out(554),
            data_im_in(43) => mul_im_out(555),
            data_im_in(44) => mul_im_out(556),
            data_im_in(45) => mul_im_out(557),
            data_im_in(46) => mul_im_out(558),
            data_im_in(47) => mul_im_out(559),
            data_im_in(48) => mul_im_out(560),
            data_im_in(49) => mul_im_out(561),
            data_im_in(50) => mul_im_out(562),
            data_im_in(51) => mul_im_out(563),
            data_im_in(52) => mul_im_out(564),
            data_im_in(53) => mul_im_out(565),
            data_im_in(54) => mul_im_out(566),
            data_im_in(55) => mul_im_out(567),
            data_im_in(56) => mul_im_out(568),
            data_im_in(57) => mul_im_out(569),
            data_im_in(58) => mul_im_out(570),
            data_im_in(59) => mul_im_out(571),
            data_im_in(60) => mul_im_out(572),
            data_im_in(61) => mul_im_out(573),
            data_im_in(62) => mul_im_out(574),
            data_im_in(63) => mul_im_out(575),
            data_re_out(0) => data_re_out(8),
            data_re_out(1) => data_re_out(40),
            data_re_out(2) => data_re_out(72),
            data_re_out(3) => data_re_out(104),
            data_re_out(4) => data_re_out(136),
            data_re_out(5) => data_re_out(168),
            data_re_out(6) => data_re_out(200),
            data_re_out(7) => data_re_out(232),
            data_re_out(8) => data_re_out(264),
            data_re_out(9) => data_re_out(296),
            data_re_out(10) => data_re_out(328),
            data_re_out(11) => data_re_out(360),
            data_re_out(12) => data_re_out(392),
            data_re_out(13) => data_re_out(424),
            data_re_out(14) => data_re_out(456),
            data_re_out(15) => data_re_out(488),
            data_re_out(16) => data_re_out(520),
            data_re_out(17) => data_re_out(552),
            data_re_out(18) => data_re_out(584),
            data_re_out(19) => data_re_out(616),
            data_re_out(20) => data_re_out(648),
            data_re_out(21) => data_re_out(680),
            data_re_out(22) => data_re_out(712),
            data_re_out(23) => data_re_out(744),
            data_re_out(24) => data_re_out(776),
            data_re_out(25) => data_re_out(808),
            data_re_out(26) => data_re_out(840),
            data_re_out(27) => data_re_out(872),
            data_re_out(28) => data_re_out(904),
            data_re_out(29) => data_re_out(936),
            data_re_out(30) => data_re_out(968),
            data_re_out(31) => data_re_out(1000),
            data_re_out(32) => data_re_out(1032),
            data_re_out(33) => data_re_out(1064),
            data_re_out(34) => data_re_out(1096),
            data_re_out(35) => data_re_out(1128),
            data_re_out(36) => data_re_out(1160),
            data_re_out(37) => data_re_out(1192),
            data_re_out(38) => data_re_out(1224),
            data_re_out(39) => data_re_out(1256),
            data_re_out(40) => data_re_out(1288),
            data_re_out(41) => data_re_out(1320),
            data_re_out(42) => data_re_out(1352),
            data_re_out(43) => data_re_out(1384),
            data_re_out(44) => data_re_out(1416),
            data_re_out(45) => data_re_out(1448),
            data_re_out(46) => data_re_out(1480),
            data_re_out(47) => data_re_out(1512),
            data_re_out(48) => data_re_out(1544),
            data_re_out(49) => data_re_out(1576),
            data_re_out(50) => data_re_out(1608),
            data_re_out(51) => data_re_out(1640),
            data_re_out(52) => data_re_out(1672),
            data_re_out(53) => data_re_out(1704),
            data_re_out(54) => data_re_out(1736),
            data_re_out(55) => data_re_out(1768),
            data_re_out(56) => data_re_out(1800),
            data_re_out(57) => data_re_out(1832),
            data_re_out(58) => data_re_out(1864),
            data_re_out(59) => data_re_out(1896),
            data_re_out(60) => data_re_out(1928),
            data_re_out(61) => data_re_out(1960),
            data_re_out(62) => data_re_out(1992),
            data_re_out(63) => data_re_out(2024),
            data_im_out(0) => data_im_out(8),
            data_im_out(1) => data_im_out(40),
            data_im_out(2) => data_im_out(72),
            data_im_out(3) => data_im_out(104),
            data_im_out(4) => data_im_out(136),
            data_im_out(5) => data_im_out(168),
            data_im_out(6) => data_im_out(200),
            data_im_out(7) => data_im_out(232),
            data_im_out(8) => data_im_out(264),
            data_im_out(9) => data_im_out(296),
            data_im_out(10) => data_im_out(328),
            data_im_out(11) => data_im_out(360),
            data_im_out(12) => data_im_out(392),
            data_im_out(13) => data_im_out(424),
            data_im_out(14) => data_im_out(456),
            data_im_out(15) => data_im_out(488),
            data_im_out(16) => data_im_out(520),
            data_im_out(17) => data_im_out(552),
            data_im_out(18) => data_im_out(584),
            data_im_out(19) => data_im_out(616),
            data_im_out(20) => data_im_out(648),
            data_im_out(21) => data_im_out(680),
            data_im_out(22) => data_im_out(712),
            data_im_out(23) => data_im_out(744),
            data_im_out(24) => data_im_out(776),
            data_im_out(25) => data_im_out(808),
            data_im_out(26) => data_im_out(840),
            data_im_out(27) => data_im_out(872),
            data_im_out(28) => data_im_out(904),
            data_im_out(29) => data_im_out(936),
            data_im_out(30) => data_im_out(968),
            data_im_out(31) => data_im_out(1000),
            data_im_out(32) => data_im_out(1032),
            data_im_out(33) => data_im_out(1064),
            data_im_out(34) => data_im_out(1096),
            data_im_out(35) => data_im_out(1128),
            data_im_out(36) => data_im_out(1160),
            data_im_out(37) => data_im_out(1192),
            data_im_out(38) => data_im_out(1224),
            data_im_out(39) => data_im_out(1256),
            data_im_out(40) => data_im_out(1288),
            data_im_out(41) => data_im_out(1320),
            data_im_out(42) => data_im_out(1352),
            data_im_out(43) => data_im_out(1384),
            data_im_out(44) => data_im_out(1416),
            data_im_out(45) => data_im_out(1448),
            data_im_out(46) => data_im_out(1480),
            data_im_out(47) => data_im_out(1512),
            data_im_out(48) => data_im_out(1544),
            data_im_out(49) => data_im_out(1576),
            data_im_out(50) => data_im_out(1608),
            data_im_out(51) => data_im_out(1640),
            data_im_out(52) => data_im_out(1672),
            data_im_out(53) => data_im_out(1704),
            data_im_out(54) => data_im_out(1736),
            data_im_out(55) => data_im_out(1768),
            data_im_out(56) => data_im_out(1800),
            data_im_out(57) => data_im_out(1832),
            data_im_out(58) => data_im_out(1864),
            data_im_out(59) => data_im_out(1896),
            data_im_out(60) => data_im_out(1928),
            data_im_out(61) => data_im_out(1960),
            data_im_out(62) => data_im_out(1992),
            data_im_out(63) => data_im_out(2024)
        );           

    URFFT_PT64_9 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(576),
            data_re_in(1) => mul_re_out(577),
            data_re_in(2) => mul_re_out(578),
            data_re_in(3) => mul_re_out(579),
            data_re_in(4) => mul_re_out(580),
            data_re_in(5) => mul_re_out(581),
            data_re_in(6) => mul_re_out(582),
            data_re_in(7) => mul_re_out(583),
            data_re_in(8) => mul_re_out(584),
            data_re_in(9) => mul_re_out(585),
            data_re_in(10) => mul_re_out(586),
            data_re_in(11) => mul_re_out(587),
            data_re_in(12) => mul_re_out(588),
            data_re_in(13) => mul_re_out(589),
            data_re_in(14) => mul_re_out(590),
            data_re_in(15) => mul_re_out(591),
            data_re_in(16) => mul_re_out(592),
            data_re_in(17) => mul_re_out(593),
            data_re_in(18) => mul_re_out(594),
            data_re_in(19) => mul_re_out(595),
            data_re_in(20) => mul_re_out(596),
            data_re_in(21) => mul_re_out(597),
            data_re_in(22) => mul_re_out(598),
            data_re_in(23) => mul_re_out(599),
            data_re_in(24) => mul_re_out(600),
            data_re_in(25) => mul_re_out(601),
            data_re_in(26) => mul_re_out(602),
            data_re_in(27) => mul_re_out(603),
            data_re_in(28) => mul_re_out(604),
            data_re_in(29) => mul_re_out(605),
            data_re_in(30) => mul_re_out(606),
            data_re_in(31) => mul_re_out(607),
            data_re_in(32) => mul_re_out(608),
            data_re_in(33) => mul_re_out(609),
            data_re_in(34) => mul_re_out(610),
            data_re_in(35) => mul_re_out(611),
            data_re_in(36) => mul_re_out(612),
            data_re_in(37) => mul_re_out(613),
            data_re_in(38) => mul_re_out(614),
            data_re_in(39) => mul_re_out(615),
            data_re_in(40) => mul_re_out(616),
            data_re_in(41) => mul_re_out(617),
            data_re_in(42) => mul_re_out(618),
            data_re_in(43) => mul_re_out(619),
            data_re_in(44) => mul_re_out(620),
            data_re_in(45) => mul_re_out(621),
            data_re_in(46) => mul_re_out(622),
            data_re_in(47) => mul_re_out(623),
            data_re_in(48) => mul_re_out(624),
            data_re_in(49) => mul_re_out(625),
            data_re_in(50) => mul_re_out(626),
            data_re_in(51) => mul_re_out(627),
            data_re_in(52) => mul_re_out(628),
            data_re_in(53) => mul_re_out(629),
            data_re_in(54) => mul_re_out(630),
            data_re_in(55) => mul_re_out(631),
            data_re_in(56) => mul_re_out(632),
            data_re_in(57) => mul_re_out(633),
            data_re_in(58) => mul_re_out(634),
            data_re_in(59) => mul_re_out(635),
            data_re_in(60) => mul_re_out(636),
            data_re_in(61) => mul_re_out(637),
            data_re_in(62) => mul_re_out(638),
            data_re_in(63) => mul_re_out(639),
            data_im_in(0) => mul_im_out(576),
            data_im_in(1) => mul_im_out(577),
            data_im_in(2) => mul_im_out(578),
            data_im_in(3) => mul_im_out(579),
            data_im_in(4) => mul_im_out(580),
            data_im_in(5) => mul_im_out(581),
            data_im_in(6) => mul_im_out(582),
            data_im_in(7) => mul_im_out(583),
            data_im_in(8) => mul_im_out(584),
            data_im_in(9) => mul_im_out(585),
            data_im_in(10) => mul_im_out(586),
            data_im_in(11) => mul_im_out(587),
            data_im_in(12) => mul_im_out(588),
            data_im_in(13) => mul_im_out(589),
            data_im_in(14) => mul_im_out(590),
            data_im_in(15) => mul_im_out(591),
            data_im_in(16) => mul_im_out(592),
            data_im_in(17) => mul_im_out(593),
            data_im_in(18) => mul_im_out(594),
            data_im_in(19) => mul_im_out(595),
            data_im_in(20) => mul_im_out(596),
            data_im_in(21) => mul_im_out(597),
            data_im_in(22) => mul_im_out(598),
            data_im_in(23) => mul_im_out(599),
            data_im_in(24) => mul_im_out(600),
            data_im_in(25) => mul_im_out(601),
            data_im_in(26) => mul_im_out(602),
            data_im_in(27) => mul_im_out(603),
            data_im_in(28) => mul_im_out(604),
            data_im_in(29) => mul_im_out(605),
            data_im_in(30) => mul_im_out(606),
            data_im_in(31) => mul_im_out(607),
            data_im_in(32) => mul_im_out(608),
            data_im_in(33) => mul_im_out(609),
            data_im_in(34) => mul_im_out(610),
            data_im_in(35) => mul_im_out(611),
            data_im_in(36) => mul_im_out(612),
            data_im_in(37) => mul_im_out(613),
            data_im_in(38) => mul_im_out(614),
            data_im_in(39) => mul_im_out(615),
            data_im_in(40) => mul_im_out(616),
            data_im_in(41) => mul_im_out(617),
            data_im_in(42) => mul_im_out(618),
            data_im_in(43) => mul_im_out(619),
            data_im_in(44) => mul_im_out(620),
            data_im_in(45) => mul_im_out(621),
            data_im_in(46) => mul_im_out(622),
            data_im_in(47) => mul_im_out(623),
            data_im_in(48) => mul_im_out(624),
            data_im_in(49) => mul_im_out(625),
            data_im_in(50) => mul_im_out(626),
            data_im_in(51) => mul_im_out(627),
            data_im_in(52) => mul_im_out(628),
            data_im_in(53) => mul_im_out(629),
            data_im_in(54) => mul_im_out(630),
            data_im_in(55) => mul_im_out(631),
            data_im_in(56) => mul_im_out(632),
            data_im_in(57) => mul_im_out(633),
            data_im_in(58) => mul_im_out(634),
            data_im_in(59) => mul_im_out(635),
            data_im_in(60) => mul_im_out(636),
            data_im_in(61) => mul_im_out(637),
            data_im_in(62) => mul_im_out(638),
            data_im_in(63) => mul_im_out(639),
            data_re_out(0) => data_re_out(9),
            data_re_out(1) => data_re_out(41),
            data_re_out(2) => data_re_out(73),
            data_re_out(3) => data_re_out(105),
            data_re_out(4) => data_re_out(137),
            data_re_out(5) => data_re_out(169),
            data_re_out(6) => data_re_out(201),
            data_re_out(7) => data_re_out(233),
            data_re_out(8) => data_re_out(265),
            data_re_out(9) => data_re_out(297),
            data_re_out(10) => data_re_out(329),
            data_re_out(11) => data_re_out(361),
            data_re_out(12) => data_re_out(393),
            data_re_out(13) => data_re_out(425),
            data_re_out(14) => data_re_out(457),
            data_re_out(15) => data_re_out(489),
            data_re_out(16) => data_re_out(521),
            data_re_out(17) => data_re_out(553),
            data_re_out(18) => data_re_out(585),
            data_re_out(19) => data_re_out(617),
            data_re_out(20) => data_re_out(649),
            data_re_out(21) => data_re_out(681),
            data_re_out(22) => data_re_out(713),
            data_re_out(23) => data_re_out(745),
            data_re_out(24) => data_re_out(777),
            data_re_out(25) => data_re_out(809),
            data_re_out(26) => data_re_out(841),
            data_re_out(27) => data_re_out(873),
            data_re_out(28) => data_re_out(905),
            data_re_out(29) => data_re_out(937),
            data_re_out(30) => data_re_out(969),
            data_re_out(31) => data_re_out(1001),
            data_re_out(32) => data_re_out(1033),
            data_re_out(33) => data_re_out(1065),
            data_re_out(34) => data_re_out(1097),
            data_re_out(35) => data_re_out(1129),
            data_re_out(36) => data_re_out(1161),
            data_re_out(37) => data_re_out(1193),
            data_re_out(38) => data_re_out(1225),
            data_re_out(39) => data_re_out(1257),
            data_re_out(40) => data_re_out(1289),
            data_re_out(41) => data_re_out(1321),
            data_re_out(42) => data_re_out(1353),
            data_re_out(43) => data_re_out(1385),
            data_re_out(44) => data_re_out(1417),
            data_re_out(45) => data_re_out(1449),
            data_re_out(46) => data_re_out(1481),
            data_re_out(47) => data_re_out(1513),
            data_re_out(48) => data_re_out(1545),
            data_re_out(49) => data_re_out(1577),
            data_re_out(50) => data_re_out(1609),
            data_re_out(51) => data_re_out(1641),
            data_re_out(52) => data_re_out(1673),
            data_re_out(53) => data_re_out(1705),
            data_re_out(54) => data_re_out(1737),
            data_re_out(55) => data_re_out(1769),
            data_re_out(56) => data_re_out(1801),
            data_re_out(57) => data_re_out(1833),
            data_re_out(58) => data_re_out(1865),
            data_re_out(59) => data_re_out(1897),
            data_re_out(60) => data_re_out(1929),
            data_re_out(61) => data_re_out(1961),
            data_re_out(62) => data_re_out(1993),
            data_re_out(63) => data_re_out(2025),
            data_im_out(0) => data_im_out(9),
            data_im_out(1) => data_im_out(41),
            data_im_out(2) => data_im_out(73),
            data_im_out(3) => data_im_out(105),
            data_im_out(4) => data_im_out(137),
            data_im_out(5) => data_im_out(169),
            data_im_out(6) => data_im_out(201),
            data_im_out(7) => data_im_out(233),
            data_im_out(8) => data_im_out(265),
            data_im_out(9) => data_im_out(297),
            data_im_out(10) => data_im_out(329),
            data_im_out(11) => data_im_out(361),
            data_im_out(12) => data_im_out(393),
            data_im_out(13) => data_im_out(425),
            data_im_out(14) => data_im_out(457),
            data_im_out(15) => data_im_out(489),
            data_im_out(16) => data_im_out(521),
            data_im_out(17) => data_im_out(553),
            data_im_out(18) => data_im_out(585),
            data_im_out(19) => data_im_out(617),
            data_im_out(20) => data_im_out(649),
            data_im_out(21) => data_im_out(681),
            data_im_out(22) => data_im_out(713),
            data_im_out(23) => data_im_out(745),
            data_im_out(24) => data_im_out(777),
            data_im_out(25) => data_im_out(809),
            data_im_out(26) => data_im_out(841),
            data_im_out(27) => data_im_out(873),
            data_im_out(28) => data_im_out(905),
            data_im_out(29) => data_im_out(937),
            data_im_out(30) => data_im_out(969),
            data_im_out(31) => data_im_out(1001),
            data_im_out(32) => data_im_out(1033),
            data_im_out(33) => data_im_out(1065),
            data_im_out(34) => data_im_out(1097),
            data_im_out(35) => data_im_out(1129),
            data_im_out(36) => data_im_out(1161),
            data_im_out(37) => data_im_out(1193),
            data_im_out(38) => data_im_out(1225),
            data_im_out(39) => data_im_out(1257),
            data_im_out(40) => data_im_out(1289),
            data_im_out(41) => data_im_out(1321),
            data_im_out(42) => data_im_out(1353),
            data_im_out(43) => data_im_out(1385),
            data_im_out(44) => data_im_out(1417),
            data_im_out(45) => data_im_out(1449),
            data_im_out(46) => data_im_out(1481),
            data_im_out(47) => data_im_out(1513),
            data_im_out(48) => data_im_out(1545),
            data_im_out(49) => data_im_out(1577),
            data_im_out(50) => data_im_out(1609),
            data_im_out(51) => data_im_out(1641),
            data_im_out(52) => data_im_out(1673),
            data_im_out(53) => data_im_out(1705),
            data_im_out(54) => data_im_out(1737),
            data_im_out(55) => data_im_out(1769),
            data_im_out(56) => data_im_out(1801),
            data_im_out(57) => data_im_out(1833),
            data_im_out(58) => data_im_out(1865),
            data_im_out(59) => data_im_out(1897),
            data_im_out(60) => data_im_out(1929),
            data_im_out(61) => data_im_out(1961),
            data_im_out(62) => data_im_out(1993),
            data_im_out(63) => data_im_out(2025)
        );           

    URFFT_PT64_10 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(640),
            data_re_in(1) => mul_re_out(641),
            data_re_in(2) => mul_re_out(642),
            data_re_in(3) => mul_re_out(643),
            data_re_in(4) => mul_re_out(644),
            data_re_in(5) => mul_re_out(645),
            data_re_in(6) => mul_re_out(646),
            data_re_in(7) => mul_re_out(647),
            data_re_in(8) => mul_re_out(648),
            data_re_in(9) => mul_re_out(649),
            data_re_in(10) => mul_re_out(650),
            data_re_in(11) => mul_re_out(651),
            data_re_in(12) => mul_re_out(652),
            data_re_in(13) => mul_re_out(653),
            data_re_in(14) => mul_re_out(654),
            data_re_in(15) => mul_re_out(655),
            data_re_in(16) => mul_re_out(656),
            data_re_in(17) => mul_re_out(657),
            data_re_in(18) => mul_re_out(658),
            data_re_in(19) => mul_re_out(659),
            data_re_in(20) => mul_re_out(660),
            data_re_in(21) => mul_re_out(661),
            data_re_in(22) => mul_re_out(662),
            data_re_in(23) => mul_re_out(663),
            data_re_in(24) => mul_re_out(664),
            data_re_in(25) => mul_re_out(665),
            data_re_in(26) => mul_re_out(666),
            data_re_in(27) => mul_re_out(667),
            data_re_in(28) => mul_re_out(668),
            data_re_in(29) => mul_re_out(669),
            data_re_in(30) => mul_re_out(670),
            data_re_in(31) => mul_re_out(671),
            data_re_in(32) => mul_re_out(672),
            data_re_in(33) => mul_re_out(673),
            data_re_in(34) => mul_re_out(674),
            data_re_in(35) => mul_re_out(675),
            data_re_in(36) => mul_re_out(676),
            data_re_in(37) => mul_re_out(677),
            data_re_in(38) => mul_re_out(678),
            data_re_in(39) => mul_re_out(679),
            data_re_in(40) => mul_re_out(680),
            data_re_in(41) => mul_re_out(681),
            data_re_in(42) => mul_re_out(682),
            data_re_in(43) => mul_re_out(683),
            data_re_in(44) => mul_re_out(684),
            data_re_in(45) => mul_re_out(685),
            data_re_in(46) => mul_re_out(686),
            data_re_in(47) => mul_re_out(687),
            data_re_in(48) => mul_re_out(688),
            data_re_in(49) => mul_re_out(689),
            data_re_in(50) => mul_re_out(690),
            data_re_in(51) => mul_re_out(691),
            data_re_in(52) => mul_re_out(692),
            data_re_in(53) => mul_re_out(693),
            data_re_in(54) => mul_re_out(694),
            data_re_in(55) => mul_re_out(695),
            data_re_in(56) => mul_re_out(696),
            data_re_in(57) => mul_re_out(697),
            data_re_in(58) => mul_re_out(698),
            data_re_in(59) => mul_re_out(699),
            data_re_in(60) => mul_re_out(700),
            data_re_in(61) => mul_re_out(701),
            data_re_in(62) => mul_re_out(702),
            data_re_in(63) => mul_re_out(703),
            data_im_in(0) => mul_im_out(640),
            data_im_in(1) => mul_im_out(641),
            data_im_in(2) => mul_im_out(642),
            data_im_in(3) => mul_im_out(643),
            data_im_in(4) => mul_im_out(644),
            data_im_in(5) => mul_im_out(645),
            data_im_in(6) => mul_im_out(646),
            data_im_in(7) => mul_im_out(647),
            data_im_in(8) => mul_im_out(648),
            data_im_in(9) => mul_im_out(649),
            data_im_in(10) => mul_im_out(650),
            data_im_in(11) => mul_im_out(651),
            data_im_in(12) => mul_im_out(652),
            data_im_in(13) => mul_im_out(653),
            data_im_in(14) => mul_im_out(654),
            data_im_in(15) => mul_im_out(655),
            data_im_in(16) => mul_im_out(656),
            data_im_in(17) => mul_im_out(657),
            data_im_in(18) => mul_im_out(658),
            data_im_in(19) => mul_im_out(659),
            data_im_in(20) => mul_im_out(660),
            data_im_in(21) => mul_im_out(661),
            data_im_in(22) => mul_im_out(662),
            data_im_in(23) => mul_im_out(663),
            data_im_in(24) => mul_im_out(664),
            data_im_in(25) => mul_im_out(665),
            data_im_in(26) => mul_im_out(666),
            data_im_in(27) => mul_im_out(667),
            data_im_in(28) => mul_im_out(668),
            data_im_in(29) => mul_im_out(669),
            data_im_in(30) => mul_im_out(670),
            data_im_in(31) => mul_im_out(671),
            data_im_in(32) => mul_im_out(672),
            data_im_in(33) => mul_im_out(673),
            data_im_in(34) => mul_im_out(674),
            data_im_in(35) => mul_im_out(675),
            data_im_in(36) => mul_im_out(676),
            data_im_in(37) => mul_im_out(677),
            data_im_in(38) => mul_im_out(678),
            data_im_in(39) => mul_im_out(679),
            data_im_in(40) => mul_im_out(680),
            data_im_in(41) => mul_im_out(681),
            data_im_in(42) => mul_im_out(682),
            data_im_in(43) => mul_im_out(683),
            data_im_in(44) => mul_im_out(684),
            data_im_in(45) => mul_im_out(685),
            data_im_in(46) => mul_im_out(686),
            data_im_in(47) => mul_im_out(687),
            data_im_in(48) => mul_im_out(688),
            data_im_in(49) => mul_im_out(689),
            data_im_in(50) => mul_im_out(690),
            data_im_in(51) => mul_im_out(691),
            data_im_in(52) => mul_im_out(692),
            data_im_in(53) => mul_im_out(693),
            data_im_in(54) => mul_im_out(694),
            data_im_in(55) => mul_im_out(695),
            data_im_in(56) => mul_im_out(696),
            data_im_in(57) => mul_im_out(697),
            data_im_in(58) => mul_im_out(698),
            data_im_in(59) => mul_im_out(699),
            data_im_in(60) => mul_im_out(700),
            data_im_in(61) => mul_im_out(701),
            data_im_in(62) => mul_im_out(702),
            data_im_in(63) => mul_im_out(703),
            data_re_out(0) => data_re_out(10),
            data_re_out(1) => data_re_out(42),
            data_re_out(2) => data_re_out(74),
            data_re_out(3) => data_re_out(106),
            data_re_out(4) => data_re_out(138),
            data_re_out(5) => data_re_out(170),
            data_re_out(6) => data_re_out(202),
            data_re_out(7) => data_re_out(234),
            data_re_out(8) => data_re_out(266),
            data_re_out(9) => data_re_out(298),
            data_re_out(10) => data_re_out(330),
            data_re_out(11) => data_re_out(362),
            data_re_out(12) => data_re_out(394),
            data_re_out(13) => data_re_out(426),
            data_re_out(14) => data_re_out(458),
            data_re_out(15) => data_re_out(490),
            data_re_out(16) => data_re_out(522),
            data_re_out(17) => data_re_out(554),
            data_re_out(18) => data_re_out(586),
            data_re_out(19) => data_re_out(618),
            data_re_out(20) => data_re_out(650),
            data_re_out(21) => data_re_out(682),
            data_re_out(22) => data_re_out(714),
            data_re_out(23) => data_re_out(746),
            data_re_out(24) => data_re_out(778),
            data_re_out(25) => data_re_out(810),
            data_re_out(26) => data_re_out(842),
            data_re_out(27) => data_re_out(874),
            data_re_out(28) => data_re_out(906),
            data_re_out(29) => data_re_out(938),
            data_re_out(30) => data_re_out(970),
            data_re_out(31) => data_re_out(1002),
            data_re_out(32) => data_re_out(1034),
            data_re_out(33) => data_re_out(1066),
            data_re_out(34) => data_re_out(1098),
            data_re_out(35) => data_re_out(1130),
            data_re_out(36) => data_re_out(1162),
            data_re_out(37) => data_re_out(1194),
            data_re_out(38) => data_re_out(1226),
            data_re_out(39) => data_re_out(1258),
            data_re_out(40) => data_re_out(1290),
            data_re_out(41) => data_re_out(1322),
            data_re_out(42) => data_re_out(1354),
            data_re_out(43) => data_re_out(1386),
            data_re_out(44) => data_re_out(1418),
            data_re_out(45) => data_re_out(1450),
            data_re_out(46) => data_re_out(1482),
            data_re_out(47) => data_re_out(1514),
            data_re_out(48) => data_re_out(1546),
            data_re_out(49) => data_re_out(1578),
            data_re_out(50) => data_re_out(1610),
            data_re_out(51) => data_re_out(1642),
            data_re_out(52) => data_re_out(1674),
            data_re_out(53) => data_re_out(1706),
            data_re_out(54) => data_re_out(1738),
            data_re_out(55) => data_re_out(1770),
            data_re_out(56) => data_re_out(1802),
            data_re_out(57) => data_re_out(1834),
            data_re_out(58) => data_re_out(1866),
            data_re_out(59) => data_re_out(1898),
            data_re_out(60) => data_re_out(1930),
            data_re_out(61) => data_re_out(1962),
            data_re_out(62) => data_re_out(1994),
            data_re_out(63) => data_re_out(2026),
            data_im_out(0) => data_im_out(10),
            data_im_out(1) => data_im_out(42),
            data_im_out(2) => data_im_out(74),
            data_im_out(3) => data_im_out(106),
            data_im_out(4) => data_im_out(138),
            data_im_out(5) => data_im_out(170),
            data_im_out(6) => data_im_out(202),
            data_im_out(7) => data_im_out(234),
            data_im_out(8) => data_im_out(266),
            data_im_out(9) => data_im_out(298),
            data_im_out(10) => data_im_out(330),
            data_im_out(11) => data_im_out(362),
            data_im_out(12) => data_im_out(394),
            data_im_out(13) => data_im_out(426),
            data_im_out(14) => data_im_out(458),
            data_im_out(15) => data_im_out(490),
            data_im_out(16) => data_im_out(522),
            data_im_out(17) => data_im_out(554),
            data_im_out(18) => data_im_out(586),
            data_im_out(19) => data_im_out(618),
            data_im_out(20) => data_im_out(650),
            data_im_out(21) => data_im_out(682),
            data_im_out(22) => data_im_out(714),
            data_im_out(23) => data_im_out(746),
            data_im_out(24) => data_im_out(778),
            data_im_out(25) => data_im_out(810),
            data_im_out(26) => data_im_out(842),
            data_im_out(27) => data_im_out(874),
            data_im_out(28) => data_im_out(906),
            data_im_out(29) => data_im_out(938),
            data_im_out(30) => data_im_out(970),
            data_im_out(31) => data_im_out(1002),
            data_im_out(32) => data_im_out(1034),
            data_im_out(33) => data_im_out(1066),
            data_im_out(34) => data_im_out(1098),
            data_im_out(35) => data_im_out(1130),
            data_im_out(36) => data_im_out(1162),
            data_im_out(37) => data_im_out(1194),
            data_im_out(38) => data_im_out(1226),
            data_im_out(39) => data_im_out(1258),
            data_im_out(40) => data_im_out(1290),
            data_im_out(41) => data_im_out(1322),
            data_im_out(42) => data_im_out(1354),
            data_im_out(43) => data_im_out(1386),
            data_im_out(44) => data_im_out(1418),
            data_im_out(45) => data_im_out(1450),
            data_im_out(46) => data_im_out(1482),
            data_im_out(47) => data_im_out(1514),
            data_im_out(48) => data_im_out(1546),
            data_im_out(49) => data_im_out(1578),
            data_im_out(50) => data_im_out(1610),
            data_im_out(51) => data_im_out(1642),
            data_im_out(52) => data_im_out(1674),
            data_im_out(53) => data_im_out(1706),
            data_im_out(54) => data_im_out(1738),
            data_im_out(55) => data_im_out(1770),
            data_im_out(56) => data_im_out(1802),
            data_im_out(57) => data_im_out(1834),
            data_im_out(58) => data_im_out(1866),
            data_im_out(59) => data_im_out(1898),
            data_im_out(60) => data_im_out(1930),
            data_im_out(61) => data_im_out(1962),
            data_im_out(62) => data_im_out(1994),
            data_im_out(63) => data_im_out(2026)
        );           

    URFFT_PT64_11 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(704),
            data_re_in(1) => mul_re_out(705),
            data_re_in(2) => mul_re_out(706),
            data_re_in(3) => mul_re_out(707),
            data_re_in(4) => mul_re_out(708),
            data_re_in(5) => mul_re_out(709),
            data_re_in(6) => mul_re_out(710),
            data_re_in(7) => mul_re_out(711),
            data_re_in(8) => mul_re_out(712),
            data_re_in(9) => mul_re_out(713),
            data_re_in(10) => mul_re_out(714),
            data_re_in(11) => mul_re_out(715),
            data_re_in(12) => mul_re_out(716),
            data_re_in(13) => mul_re_out(717),
            data_re_in(14) => mul_re_out(718),
            data_re_in(15) => mul_re_out(719),
            data_re_in(16) => mul_re_out(720),
            data_re_in(17) => mul_re_out(721),
            data_re_in(18) => mul_re_out(722),
            data_re_in(19) => mul_re_out(723),
            data_re_in(20) => mul_re_out(724),
            data_re_in(21) => mul_re_out(725),
            data_re_in(22) => mul_re_out(726),
            data_re_in(23) => mul_re_out(727),
            data_re_in(24) => mul_re_out(728),
            data_re_in(25) => mul_re_out(729),
            data_re_in(26) => mul_re_out(730),
            data_re_in(27) => mul_re_out(731),
            data_re_in(28) => mul_re_out(732),
            data_re_in(29) => mul_re_out(733),
            data_re_in(30) => mul_re_out(734),
            data_re_in(31) => mul_re_out(735),
            data_re_in(32) => mul_re_out(736),
            data_re_in(33) => mul_re_out(737),
            data_re_in(34) => mul_re_out(738),
            data_re_in(35) => mul_re_out(739),
            data_re_in(36) => mul_re_out(740),
            data_re_in(37) => mul_re_out(741),
            data_re_in(38) => mul_re_out(742),
            data_re_in(39) => mul_re_out(743),
            data_re_in(40) => mul_re_out(744),
            data_re_in(41) => mul_re_out(745),
            data_re_in(42) => mul_re_out(746),
            data_re_in(43) => mul_re_out(747),
            data_re_in(44) => mul_re_out(748),
            data_re_in(45) => mul_re_out(749),
            data_re_in(46) => mul_re_out(750),
            data_re_in(47) => mul_re_out(751),
            data_re_in(48) => mul_re_out(752),
            data_re_in(49) => mul_re_out(753),
            data_re_in(50) => mul_re_out(754),
            data_re_in(51) => mul_re_out(755),
            data_re_in(52) => mul_re_out(756),
            data_re_in(53) => mul_re_out(757),
            data_re_in(54) => mul_re_out(758),
            data_re_in(55) => mul_re_out(759),
            data_re_in(56) => mul_re_out(760),
            data_re_in(57) => mul_re_out(761),
            data_re_in(58) => mul_re_out(762),
            data_re_in(59) => mul_re_out(763),
            data_re_in(60) => mul_re_out(764),
            data_re_in(61) => mul_re_out(765),
            data_re_in(62) => mul_re_out(766),
            data_re_in(63) => mul_re_out(767),
            data_im_in(0) => mul_im_out(704),
            data_im_in(1) => mul_im_out(705),
            data_im_in(2) => mul_im_out(706),
            data_im_in(3) => mul_im_out(707),
            data_im_in(4) => mul_im_out(708),
            data_im_in(5) => mul_im_out(709),
            data_im_in(6) => mul_im_out(710),
            data_im_in(7) => mul_im_out(711),
            data_im_in(8) => mul_im_out(712),
            data_im_in(9) => mul_im_out(713),
            data_im_in(10) => mul_im_out(714),
            data_im_in(11) => mul_im_out(715),
            data_im_in(12) => mul_im_out(716),
            data_im_in(13) => mul_im_out(717),
            data_im_in(14) => mul_im_out(718),
            data_im_in(15) => mul_im_out(719),
            data_im_in(16) => mul_im_out(720),
            data_im_in(17) => mul_im_out(721),
            data_im_in(18) => mul_im_out(722),
            data_im_in(19) => mul_im_out(723),
            data_im_in(20) => mul_im_out(724),
            data_im_in(21) => mul_im_out(725),
            data_im_in(22) => mul_im_out(726),
            data_im_in(23) => mul_im_out(727),
            data_im_in(24) => mul_im_out(728),
            data_im_in(25) => mul_im_out(729),
            data_im_in(26) => mul_im_out(730),
            data_im_in(27) => mul_im_out(731),
            data_im_in(28) => mul_im_out(732),
            data_im_in(29) => mul_im_out(733),
            data_im_in(30) => mul_im_out(734),
            data_im_in(31) => mul_im_out(735),
            data_im_in(32) => mul_im_out(736),
            data_im_in(33) => mul_im_out(737),
            data_im_in(34) => mul_im_out(738),
            data_im_in(35) => mul_im_out(739),
            data_im_in(36) => mul_im_out(740),
            data_im_in(37) => mul_im_out(741),
            data_im_in(38) => mul_im_out(742),
            data_im_in(39) => mul_im_out(743),
            data_im_in(40) => mul_im_out(744),
            data_im_in(41) => mul_im_out(745),
            data_im_in(42) => mul_im_out(746),
            data_im_in(43) => mul_im_out(747),
            data_im_in(44) => mul_im_out(748),
            data_im_in(45) => mul_im_out(749),
            data_im_in(46) => mul_im_out(750),
            data_im_in(47) => mul_im_out(751),
            data_im_in(48) => mul_im_out(752),
            data_im_in(49) => mul_im_out(753),
            data_im_in(50) => mul_im_out(754),
            data_im_in(51) => mul_im_out(755),
            data_im_in(52) => mul_im_out(756),
            data_im_in(53) => mul_im_out(757),
            data_im_in(54) => mul_im_out(758),
            data_im_in(55) => mul_im_out(759),
            data_im_in(56) => mul_im_out(760),
            data_im_in(57) => mul_im_out(761),
            data_im_in(58) => mul_im_out(762),
            data_im_in(59) => mul_im_out(763),
            data_im_in(60) => mul_im_out(764),
            data_im_in(61) => mul_im_out(765),
            data_im_in(62) => mul_im_out(766),
            data_im_in(63) => mul_im_out(767),
            data_re_out(0) => data_re_out(11),
            data_re_out(1) => data_re_out(43),
            data_re_out(2) => data_re_out(75),
            data_re_out(3) => data_re_out(107),
            data_re_out(4) => data_re_out(139),
            data_re_out(5) => data_re_out(171),
            data_re_out(6) => data_re_out(203),
            data_re_out(7) => data_re_out(235),
            data_re_out(8) => data_re_out(267),
            data_re_out(9) => data_re_out(299),
            data_re_out(10) => data_re_out(331),
            data_re_out(11) => data_re_out(363),
            data_re_out(12) => data_re_out(395),
            data_re_out(13) => data_re_out(427),
            data_re_out(14) => data_re_out(459),
            data_re_out(15) => data_re_out(491),
            data_re_out(16) => data_re_out(523),
            data_re_out(17) => data_re_out(555),
            data_re_out(18) => data_re_out(587),
            data_re_out(19) => data_re_out(619),
            data_re_out(20) => data_re_out(651),
            data_re_out(21) => data_re_out(683),
            data_re_out(22) => data_re_out(715),
            data_re_out(23) => data_re_out(747),
            data_re_out(24) => data_re_out(779),
            data_re_out(25) => data_re_out(811),
            data_re_out(26) => data_re_out(843),
            data_re_out(27) => data_re_out(875),
            data_re_out(28) => data_re_out(907),
            data_re_out(29) => data_re_out(939),
            data_re_out(30) => data_re_out(971),
            data_re_out(31) => data_re_out(1003),
            data_re_out(32) => data_re_out(1035),
            data_re_out(33) => data_re_out(1067),
            data_re_out(34) => data_re_out(1099),
            data_re_out(35) => data_re_out(1131),
            data_re_out(36) => data_re_out(1163),
            data_re_out(37) => data_re_out(1195),
            data_re_out(38) => data_re_out(1227),
            data_re_out(39) => data_re_out(1259),
            data_re_out(40) => data_re_out(1291),
            data_re_out(41) => data_re_out(1323),
            data_re_out(42) => data_re_out(1355),
            data_re_out(43) => data_re_out(1387),
            data_re_out(44) => data_re_out(1419),
            data_re_out(45) => data_re_out(1451),
            data_re_out(46) => data_re_out(1483),
            data_re_out(47) => data_re_out(1515),
            data_re_out(48) => data_re_out(1547),
            data_re_out(49) => data_re_out(1579),
            data_re_out(50) => data_re_out(1611),
            data_re_out(51) => data_re_out(1643),
            data_re_out(52) => data_re_out(1675),
            data_re_out(53) => data_re_out(1707),
            data_re_out(54) => data_re_out(1739),
            data_re_out(55) => data_re_out(1771),
            data_re_out(56) => data_re_out(1803),
            data_re_out(57) => data_re_out(1835),
            data_re_out(58) => data_re_out(1867),
            data_re_out(59) => data_re_out(1899),
            data_re_out(60) => data_re_out(1931),
            data_re_out(61) => data_re_out(1963),
            data_re_out(62) => data_re_out(1995),
            data_re_out(63) => data_re_out(2027),
            data_im_out(0) => data_im_out(11),
            data_im_out(1) => data_im_out(43),
            data_im_out(2) => data_im_out(75),
            data_im_out(3) => data_im_out(107),
            data_im_out(4) => data_im_out(139),
            data_im_out(5) => data_im_out(171),
            data_im_out(6) => data_im_out(203),
            data_im_out(7) => data_im_out(235),
            data_im_out(8) => data_im_out(267),
            data_im_out(9) => data_im_out(299),
            data_im_out(10) => data_im_out(331),
            data_im_out(11) => data_im_out(363),
            data_im_out(12) => data_im_out(395),
            data_im_out(13) => data_im_out(427),
            data_im_out(14) => data_im_out(459),
            data_im_out(15) => data_im_out(491),
            data_im_out(16) => data_im_out(523),
            data_im_out(17) => data_im_out(555),
            data_im_out(18) => data_im_out(587),
            data_im_out(19) => data_im_out(619),
            data_im_out(20) => data_im_out(651),
            data_im_out(21) => data_im_out(683),
            data_im_out(22) => data_im_out(715),
            data_im_out(23) => data_im_out(747),
            data_im_out(24) => data_im_out(779),
            data_im_out(25) => data_im_out(811),
            data_im_out(26) => data_im_out(843),
            data_im_out(27) => data_im_out(875),
            data_im_out(28) => data_im_out(907),
            data_im_out(29) => data_im_out(939),
            data_im_out(30) => data_im_out(971),
            data_im_out(31) => data_im_out(1003),
            data_im_out(32) => data_im_out(1035),
            data_im_out(33) => data_im_out(1067),
            data_im_out(34) => data_im_out(1099),
            data_im_out(35) => data_im_out(1131),
            data_im_out(36) => data_im_out(1163),
            data_im_out(37) => data_im_out(1195),
            data_im_out(38) => data_im_out(1227),
            data_im_out(39) => data_im_out(1259),
            data_im_out(40) => data_im_out(1291),
            data_im_out(41) => data_im_out(1323),
            data_im_out(42) => data_im_out(1355),
            data_im_out(43) => data_im_out(1387),
            data_im_out(44) => data_im_out(1419),
            data_im_out(45) => data_im_out(1451),
            data_im_out(46) => data_im_out(1483),
            data_im_out(47) => data_im_out(1515),
            data_im_out(48) => data_im_out(1547),
            data_im_out(49) => data_im_out(1579),
            data_im_out(50) => data_im_out(1611),
            data_im_out(51) => data_im_out(1643),
            data_im_out(52) => data_im_out(1675),
            data_im_out(53) => data_im_out(1707),
            data_im_out(54) => data_im_out(1739),
            data_im_out(55) => data_im_out(1771),
            data_im_out(56) => data_im_out(1803),
            data_im_out(57) => data_im_out(1835),
            data_im_out(58) => data_im_out(1867),
            data_im_out(59) => data_im_out(1899),
            data_im_out(60) => data_im_out(1931),
            data_im_out(61) => data_im_out(1963),
            data_im_out(62) => data_im_out(1995),
            data_im_out(63) => data_im_out(2027)
        );           

    URFFT_PT64_12 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(768),
            data_re_in(1) => mul_re_out(769),
            data_re_in(2) => mul_re_out(770),
            data_re_in(3) => mul_re_out(771),
            data_re_in(4) => mul_re_out(772),
            data_re_in(5) => mul_re_out(773),
            data_re_in(6) => mul_re_out(774),
            data_re_in(7) => mul_re_out(775),
            data_re_in(8) => mul_re_out(776),
            data_re_in(9) => mul_re_out(777),
            data_re_in(10) => mul_re_out(778),
            data_re_in(11) => mul_re_out(779),
            data_re_in(12) => mul_re_out(780),
            data_re_in(13) => mul_re_out(781),
            data_re_in(14) => mul_re_out(782),
            data_re_in(15) => mul_re_out(783),
            data_re_in(16) => mul_re_out(784),
            data_re_in(17) => mul_re_out(785),
            data_re_in(18) => mul_re_out(786),
            data_re_in(19) => mul_re_out(787),
            data_re_in(20) => mul_re_out(788),
            data_re_in(21) => mul_re_out(789),
            data_re_in(22) => mul_re_out(790),
            data_re_in(23) => mul_re_out(791),
            data_re_in(24) => mul_re_out(792),
            data_re_in(25) => mul_re_out(793),
            data_re_in(26) => mul_re_out(794),
            data_re_in(27) => mul_re_out(795),
            data_re_in(28) => mul_re_out(796),
            data_re_in(29) => mul_re_out(797),
            data_re_in(30) => mul_re_out(798),
            data_re_in(31) => mul_re_out(799),
            data_re_in(32) => mul_re_out(800),
            data_re_in(33) => mul_re_out(801),
            data_re_in(34) => mul_re_out(802),
            data_re_in(35) => mul_re_out(803),
            data_re_in(36) => mul_re_out(804),
            data_re_in(37) => mul_re_out(805),
            data_re_in(38) => mul_re_out(806),
            data_re_in(39) => mul_re_out(807),
            data_re_in(40) => mul_re_out(808),
            data_re_in(41) => mul_re_out(809),
            data_re_in(42) => mul_re_out(810),
            data_re_in(43) => mul_re_out(811),
            data_re_in(44) => mul_re_out(812),
            data_re_in(45) => mul_re_out(813),
            data_re_in(46) => mul_re_out(814),
            data_re_in(47) => mul_re_out(815),
            data_re_in(48) => mul_re_out(816),
            data_re_in(49) => mul_re_out(817),
            data_re_in(50) => mul_re_out(818),
            data_re_in(51) => mul_re_out(819),
            data_re_in(52) => mul_re_out(820),
            data_re_in(53) => mul_re_out(821),
            data_re_in(54) => mul_re_out(822),
            data_re_in(55) => mul_re_out(823),
            data_re_in(56) => mul_re_out(824),
            data_re_in(57) => mul_re_out(825),
            data_re_in(58) => mul_re_out(826),
            data_re_in(59) => mul_re_out(827),
            data_re_in(60) => mul_re_out(828),
            data_re_in(61) => mul_re_out(829),
            data_re_in(62) => mul_re_out(830),
            data_re_in(63) => mul_re_out(831),
            data_im_in(0) => mul_im_out(768),
            data_im_in(1) => mul_im_out(769),
            data_im_in(2) => mul_im_out(770),
            data_im_in(3) => mul_im_out(771),
            data_im_in(4) => mul_im_out(772),
            data_im_in(5) => mul_im_out(773),
            data_im_in(6) => mul_im_out(774),
            data_im_in(7) => mul_im_out(775),
            data_im_in(8) => mul_im_out(776),
            data_im_in(9) => mul_im_out(777),
            data_im_in(10) => mul_im_out(778),
            data_im_in(11) => mul_im_out(779),
            data_im_in(12) => mul_im_out(780),
            data_im_in(13) => mul_im_out(781),
            data_im_in(14) => mul_im_out(782),
            data_im_in(15) => mul_im_out(783),
            data_im_in(16) => mul_im_out(784),
            data_im_in(17) => mul_im_out(785),
            data_im_in(18) => mul_im_out(786),
            data_im_in(19) => mul_im_out(787),
            data_im_in(20) => mul_im_out(788),
            data_im_in(21) => mul_im_out(789),
            data_im_in(22) => mul_im_out(790),
            data_im_in(23) => mul_im_out(791),
            data_im_in(24) => mul_im_out(792),
            data_im_in(25) => mul_im_out(793),
            data_im_in(26) => mul_im_out(794),
            data_im_in(27) => mul_im_out(795),
            data_im_in(28) => mul_im_out(796),
            data_im_in(29) => mul_im_out(797),
            data_im_in(30) => mul_im_out(798),
            data_im_in(31) => mul_im_out(799),
            data_im_in(32) => mul_im_out(800),
            data_im_in(33) => mul_im_out(801),
            data_im_in(34) => mul_im_out(802),
            data_im_in(35) => mul_im_out(803),
            data_im_in(36) => mul_im_out(804),
            data_im_in(37) => mul_im_out(805),
            data_im_in(38) => mul_im_out(806),
            data_im_in(39) => mul_im_out(807),
            data_im_in(40) => mul_im_out(808),
            data_im_in(41) => mul_im_out(809),
            data_im_in(42) => mul_im_out(810),
            data_im_in(43) => mul_im_out(811),
            data_im_in(44) => mul_im_out(812),
            data_im_in(45) => mul_im_out(813),
            data_im_in(46) => mul_im_out(814),
            data_im_in(47) => mul_im_out(815),
            data_im_in(48) => mul_im_out(816),
            data_im_in(49) => mul_im_out(817),
            data_im_in(50) => mul_im_out(818),
            data_im_in(51) => mul_im_out(819),
            data_im_in(52) => mul_im_out(820),
            data_im_in(53) => mul_im_out(821),
            data_im_in(54) => mul_im_out(822),
            data_im_in(55) => mul_im_out(823),
            data_im_in(56) => mul_im_out(824),
            data_im_in(57) => mul_im_out(825),
            data_im_in(58) => mul_im_out(826),
            data_im_in(59) => mul_im_out(827),
            data_im_in(60) => mul_im_out(828),
            data_im_in(61) => mul_im_out(829),
            data_im_in(62) => mul_im_out(830),
            data_im_in(63) => mul_im_out(831),
            data_re_out(0) => data_re_out(12),
            data_re_out(1) => data_re_out(44),
            data_re_out(2) => data_re_out(76),
            data_re_out(3) => data_re_out(108),
            data_re_out(4) => data_re_out(140),
            data_re_out(5) => data_re_out(172),
            data_re_out(6) => data_re_out(204),
            data_re_out(7) => data_re_out(236),
            data_re_out(8) => data_re_out(268),
            data_re_out(9) => data_re_out(300),
            data_re_out(10) => data_re_out(332),
            data_re_out(11) => data_re_out(364),
            data_re_out(12) => data_re_out(396),
            data_re_out(13) => data_re_out(428),
            data_re_out(14) => data_re_out(460),
            data_re_out(15) => data_re_out(492),
            data_re_out(16) => data_re_out(524),
            data_re_out(17) => data_re_out(556),
            data_re_out(18) => data_re_out(588),
            data_re_out(19) => data_re_out(620),
            data_re_out(20) => data_re_out(652),
            data_re_out(21) => data_re_out(684),
            data_re_out(22) => data_re_out(716),
            data_re_out(23) => data_re_out(748),
            data_re_out(24) => data_re_out(780),
            data_re_out(25) => data_re_out(812),
            data_re_out(26) => data_re_out(844),
            data_re_out(27) => data_re_out(876),
            data_re_out(28) => data_re_out(908),
            data_re_out(29) => data_re_out(940),
            data_re_out(30) => data_re_out(972),
            data_re_out(31) => data_re_out(1004),
            data_re_out(32) => data_re_out(1036),
            data_re_out(33) => data_re_out(1068),
            data_re_out(34) => data_re_out(1100),
            data_re_out(35) => data_re_out(1132),
            data_re_out(36) => data_re_out(1164),
            data_re_out(37) => data_re_out(1196),
            data_re_out(38) => data_re_out(1228),
            data_re_out(39) => data_re_out(1260),
            data_re_out(40) => data_re_out(1292),
            data_re_out(41) => data_re_out(1324),
            data_re_out(42) => data_re_out(1356),
            data_re_out(43) => data_re_out(1388),
            data_re_out(44) => data_re_out(1420),
            data_re_out(45) => data_re_out(1452),
            data_re_out(46) => data_re_out(1484),
            data_re_out(47) => data_re_out(1516),
            data_re_out(48) => data_re_out(1548),
            data_re_out(49) => data_re_out(1580),
            data_re_out(50) => data_re_out(1612),
            data_re_out(51) => data_re_out(1644),
            data_re_out(52) => data_re_out(1676),
            data_re_out(53) => data_re_out(1708),
            data_re_out(54) => data_re_out(1740),
            data_re_out(55) => data_re_out(1772),
            data_re_out(56) => data_re_out(1804),
            data_re_out(57) => data_re_out(1836),
            data_re_out(58) => data_re_out(1868),
            data_re_out(59) => data_re_out(1900),
            data_re_out(60) => data_re_out(1932),
            data_re_out(61) => data_re_out(1964),
            data_re_out(62) => data_re_out(1996),
            data_re_out(63) => data_re_out(2028),
            data_im_out(0) => data_im_out(12),
            data_im_out(1) => data_im_out(44),
            data_im_out(2) => data_im_out(76),
            data_im_out(3) => data_im_out(108),
            data_im_out(4) => data_im_out(140),
            data_im_out(5) => data_im_out(172),
            data_im_out(6) => data_im_out(204),
            data_im_out(7) => data_im_out(236),
            data_im_out(8) => data_im_out(268),
            data_im_out(9) => data_im_out(300),
            data_im_out(10) => data_im_out(332),
            data_im_out(11) => data_im_out(364),
            data_im_out(12) => data_im_out(396),
            data_im_out(13) => data_im_out(428),
            data_im_out(14) => data_im_out(460),
            data_im_out(15) => data_im_out(492),
            data_im_out(16) => data_im_out(524),
            data_im_out(17) => data_im_out(556),
            data_im_out(18) => data_im_out(588),
            data_im_out(19) => data_im_out(620),
            data_im_out(20) => data_im_out(652),
            data_im_out(21) => data_im_out(684),
            data_im_out(22) => data_im_out(716),
            data_im_out(23) => data_im_out(748),
            data_im_out(24) => data_im_out(780),
            data_im_out(25) => data_im_out(812),
            data_im_out(26) => data_im_out(844),
            data_im_out(27) => data_im_out(876),
            data_im_out(28) => data_im_out(908),
            data_im_out(29) => data_im_out(940),
            data_im_out(30) => data_im_out(972),
            data_im_out(31) => data_im_out(1004),
            data_im_out(32) => data_im_out(1036),
            data_im_out(33) => data_im_out(1068),
            data_im_out(34) => data_im_out(1100),
            data_im_out(35) => data_im_out(1132),
            data_im_out(36) => data_im_out(1164),
            data_im_out(37) => data_im_out(1196),
            data_im_out(38) => data_im_out(1228),
            data_im_out(39) => data_im_out(1260),
            data_im_out(40) => data_im_out(1292),
            data_im_out(41) => data_im_out(1324),
            data_im_out(42) => data_im_out(1356),
            data_im_out(43) => data_im_out(1388),
            data_im_out(44) => data_im_out(1420),
            data_im_out(45) => data_im_out(1452),
            data_im_out(46) => data_im_out(1484),
            data_im_out(47) => data_im_out(1516),
            data_im_out(48) => data_im_out(1548),
            data_im_out(49) => data_im_out(1580),
            data_im_out(50) => data_im_out(1612),
            data_im_out(51) => data_im_out(1644),
            data_im_out(52) => data_im_out(1676),
            data_im_out(53) => data_im_out(1708),
            data_im_out(54) => data_im_out(1740),
            data_im_out(55) => data_im_out(1772),
            data_im_out(56) => data_im_out(1804),
            data_im_out(57) => data_im_out(1836),
            data_im_out(58) => data_im_out(1868),
            data_im_out(59) => data_im_out(1900),
            data_im_out(60) => data_im_out(1932),
            data_im_out(61) => data_im_out(1964),
            data_im_out(62) => data_im_out(1996),
            data_im_out(63) => data_im_out(2028)
        );           

    URFFT_PT64_13 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(832),
            data_re_in(1) => mul_re_out(833),
            data_re_in(2) => mul_re_out(834),
            data_re_in(3) => mul_re_out(835),
            data_re_in(4) => mul_re_out(836),
            data_re_in(5) => mul_re_out(837),
            data_re_in(6) => mul_re_out(838),
            data_re_in(7) => mul_re_out(839),
            data_re_in(8) => mul_re_out(840),
            data_re_in(9) => mul_re_out(841),
            data_re_in(10) => mul_re_out(842),
            data_re_in(11) => mul_re_out(843),
            data_re_in(12) => mul_re_out(844),
            data_re_in(13) => mul_re_out(845),
            data_re_in(14) => mul_re_out(846),
            data_re_in(15) => mul_re_out(847),
            data_re_in(16) => mul_re_out(848),
            data_re_in(17) => mul_re_out(849),
            data_re_in(18) => mul_re_out(850),
            data_re_in(19) => mul_re_out(851),
            data_re_in(20) => mul_re_out(852),
            data_re_in(21) => mul_re_out(853),
            data_re_in(22) => mul_re_out(854),
            data_re_in(23) => mul_re_out(855),
            data_re_in(24) => mul_re_out(856),
            data_re_in(25) => mul_re_out(857),
            data_re_in(26) => mul_re_out(858),
            data_re_in(27) => mul_re_out(859),
            data_re_in(28) => mul_re_out(860),
            data_re_in(29) => mul_re_out(861),
            data_re_in(30) => mul_re_out(862),
            data_re_in(31) => mul_re_out(863),
            data_re_in(32) => mul_re_out(864),
            data_re_in(33) => mul_re_out(865),
            data_re_in(34) => mul_re_out(866),
            data_re_in(35) => mul_re_out(867),
            data_re_in(36) => mul_re_out(868),
            data_re_in(37) => mul_re_out(869),
            data_re_in(38) => mul_re_out(870),
            data_re_in(39) => mul_re_out(871),
            data_re_in(40) => mul_re_out(872),
            data_re_in(41) => mul_re_out(873),
            data_re_in(42) => mul_re_out(874),
            data_re_in(43) => mul_re_out(875),
            data_re_in(44) => mul_re_out(876),
            data_re_in(45) => mul_re_out(877),
            data_re_in(46) => mul_re_out(878),
            data_re_in(47) => mul_re_out(879),
            data_re_in(48) => mul_re_out(880),
            data_re_in(49) => mul_re_out(881),
            data_re_in(50) => mul_re_out(882),
            data_re_in(51) => mul_re_out(883),
            data_re_in(52) => mul_re_out(884),
            data_re_in(53) => mul_re_out(885),
            data_re_in(54) => mul_re_out(886),
            data_re_in(55) => mul_re_out(887),
            data_re_in(56) => mul_re_out(888),
            data_re_in(57) => mul_re_out(889),
            data_re_in(58) => mul_re_out(890),
            data_re_in(59) => mul_re_out(891),
            data_re_in(60) => mul_re_out(892),
            data_re_in(61) => mul_re_out(893),
            data_re_in(62) => mul_re_out(894),
            data_re_in(63) => mul_re_out(895),
            data_im_in(0) => mul_im_out(832),
            data_im_in(1) => mul_im_out(833),
            data_im_in(2) => mul_im_out(834),
            data_im_in(3) => mul_im_out(835),
            data_im_in(4) => mul_im_out(836),
            data_im_in(5) => mul_im_out(837),
            data_im_in(6) => mul_im_out(838),
            data_im_in(7) => mul_im_out(839),
            data_im_in(8) => mul_im_out(840),
            data_im_in(9) => mul_im_out(841),
            data_im_in(10) => mul_im_out(842),
            data_im_in(11) => mul_im_out(843),
            data_im_in(12) => mul_im_out(844),
            data_im_in(13) => mul_im_out(845),
            data_im_in(14) => mul_im_out(846),
            data_im_in(15) => mul_im_out(847),
            data_im_in(16) => mul_im_out(848),
            data_im_in(17) => mul_im_out(849),
            data_im_in(18) => mul_im_out(850),
            data_im_in(19) => mul_im_out(851),
            data_im_in(20) => mul_im_out(852),
            data_im_in(21) => mul_im_out(853),
            data_im_in(22) => mul_im_out(854),
            data_im_in(23) => mul_im_out(855),
            data_im_in(24) => mul_im_out(856),
            data_im_in(25) => mul_im_out(857),
            data_im_in(26) => mul_im_out(858),
            data_im_in(27) => mul_im_out(859),
            data_im_in(28) => mul_im_out(860),
            data_im_in(29) => mul_im_out(861),
            data_im_in(30) => mul_im_out(862),
            data_im_in(31) => mul_im_out(863),
            data_im_in(32) => mul_im_out(864),
            data_im_in(33) => mul_im_out(865),
            data_im_in(34) => mul_im_out(866),
            data_im_in(35) => mul_im_out(867),
            data_im_in(36) => mul_im_out(868),
            data_im_in(37) => mul_im_out(869),
            data_im_in(38) => mul_im_out(870),
            data_im_in(39) => mul_im_out(871),
            data_im_in(40) => mul_im_out(872),
            data_im_in(41) => mul_im_out(873),
            data_im_in(42) => mul_im_out(874),
            data_im_in(43) => mul_im_out(875),
            data_im_in(44) => mul_im_out(876),
            data_im_in(45) => mul_im_out(877),
            data_im_in(46) => mul_im_out(878),
            data_im_in(47) => mul_im_out(879),
            data_im_in(48) => mul_im_out(880),
            data_im_in(49) => mul_im_out(881),
            data_im_in(50) => mul_im_out(882),
            data_im_in(51) => mul_im_out(883),
            data_im_in(52) => mul_im_out(884),
            data_im_in(53) => mul_im_out(885),
            data_im_in(54) => mul_im_out(886),
            data_im_in(55) => mul_im_out(887),
            data_im_in(56) => mul_im_out(888),
            data_im_in(57) => mul_im_out(889),
            data_im_in(58) => mul_im_out(890),
            data_im_in(59) => mul_im_out(891),
            data_im_in(60) => mul_im_out(892),
            data_im_in(61) => mul_im_out(893),
            data_im_in(62) => mul_im_out(894),
            data_im_in(63) => mul_im_out(895),
            data_re_out(0) => data_re_out(13),
            data_re_out(1) => data_re_out(45),
            data_re_out(2) => data_re_out(77),
            data_re_out(3) => data_re_out(109),
            data_re_out(4) => data_re_out(141),
            data_re_out(5) => data_re_out(173),
            data_re_out(6) => data_re_out(205),
            data_re_out(7) => data_re_out(237),
            data_re_out(8) => data_re_out(269),
            data_re_out(9) => data_re_out(301),
            data_re_out(10) => data_re_out(333),
            data_re_out(11) => data_re_out(365),
            data_re_out(12) => data_re_out(397),
            data_re_out(13) => data_re_out(429),
            data_re_out(14) => data_re_out(461),
            data_re_out(15) => data_re_out(493),
            data_re_out(16) => data_re_out(525),
            data_re_out(17) => data_re_out(557),
            data_re_out(18) => data_re_out(589),
            data_re_out(19) => data_re_out(621),
            data_re_out(20) => data_re_out(653),
            data_re_out(21) => data_re_out(685),
            data_re_out(22) => data_re_out(717),
            data_re_out(23) => data_re_out(749),
            data_re_out(24) => data_re_out(781),
            data_re_out(25) => data_re_out(813),
            data_re_out(26) => data_re_out(845),
            data_re_out(27) => data_re_out(877),
            data_re_out(28) => data_re_out(909),
            data_re_out(29) => data_re_out(941),
            data_re_out(30) => data_re_out(973),
            data_re_out(31) => data_re_out(1005),
            data_re_out(32) => data_re_out(1037),
            data_re_out(33) => data_re_out(1069),
            data_re_out(34) => data_re_out(1101),
            data_re_out(35) => data_re_out(1133),
            data_re_out(36) => data_re_out(1165),
            data_re_out(37) => data_re_out(1197),
            data_re_out(38) => data_re_out(1229),
            data_re_out(39) => data_re_out(1261),
            data_re_out(40) => data_re_out(1293),
            data_re_out(41) => data_re_out(1325),
            data_re_out(42) => data_re_out(1357),
            data_re_out(43) => data_re_out(1389),
            data_re_out(44) => data_re_out(1421),
            data_re_out(45) => data_re_out(1453),
            data_re_out(46) => data_re_out(1485),
            data_re_out(47) => data_re_out(1517),
            data_re_out(48) => data_re_out(1549),
            data_re_out(49) => data_re_out(1581),
            data_re_out(50) => data_re_out(1613),
            data_re_out(51) => data_re_out(1645),
            data_re_out(52) => data_re_out(1677),
            data_re_out(53) => data_re_out(1709),
            data_re_out(54) => data_re_out(1741),
            data_re_out(55) => data_re_out(1773),
            data_re_out(56) => data_re_out(1805),
            data_re_out(57) => data_re_out(1837),
            data_re_out(58) => data_re_out(1869),
            data_re_out(59) => data_re_out(1901),
            data_re_out(60) => data_re_out(1933),
            data_re_out(61) => data_re_out(1965),
            data_re_out(62) => data_re_out(1997),
            data_re_out(63) => data_re_out(2029),
            data_im_out(0) => data_im_out(13),
            data_im_out(1) => data_im_out(45),
            data_im_out(2) => data_im_out(77),
            data_im_out(3) => data_im_out(109),
            data_im_out(4) => data_im_out(141),
            data_im_out(5) => data_im_out(173),
            data_im_out(6) => data_im_out(205),
            data_im_out(7) => data_im_out(237),
            data_im_out(8) => data_im_out(269),
            data_im_out(9) => data_im_out(301),
            data_im_out(10) => data_im_out(333),
            data_im_out(11) => data_im_out(365),
            data_im_out(12) => data_im_out(397),
            data_im_out(13) => data_im_out(429),
            data_im_out(14) => data_im_out(461),
            data_im_out(15) => data_im_out(493),
            data_im_out(16) => data_im_out(525),
            data_im_out(17) => data_im_out(557),
            data_im_out(18) => data_im_out(589),
            data_im_out(19) => data_im_out(621),
            data_im_out(20) => data_im_out(653),
            data_im_out(21) => data_im_out(685),
            data_im_out(22) => data_im_out(717),
            data_im_out(23) => data_im_out(749),
            data_im_out(24) => data_im_out(781),
            data_im_out(25) => data_im_out(813),
            data_im_out(26) => data_im_out(845),
            data_im_out(27) => data_im_out(877),
            data_im_out(28) => data_im_out(909),
            data_im_out(29) => data_im_out(941),
            data_im_out(30) => data_im_out(973),
            data_im_out(31) => data_im_out(1005),
            data_im_out(32) => data_im_out(1037),
            data_im_out(33) => data_im_out(1069),
            data_im_out(34) => data_im_out(1101),
            data_im_out(35) => data_im_out(1133),
            data_im_out(36) => data_im_out(1165),
            data_im_out(37) => data_im_out(1197),
            data_im_out(38) => data_im_out(1229),
            data_im_out(39) => data_im_out(1261),
            data_im_out(40) => data_im_out(1293),
            data_im_out(41) => data_im_out(1325),
            data_im_out(42) => data_im_out(1357),
            data_im_out(43) => data_im_out(1389),
            data_im_out(44) => data_im_out(1421),
            data_im_out(45) => data_im_out(1453),
            data_im_out(46) => data_im_out(1485),
            data_im_out(47) => data_im_out(1517),
            data_im_out(48) => data_im_out(1549),
            data_im_out(49) => data_im_out(1581),
            data_im_out(50) => data_im_out(1613),
            data_im_out(51) => data_im_out(1645),
            data_im_out(52) => data_im_out(1677),
            data_im_out(53) => data_im_out(1709),
            data_im_out(54) => data_im_out(1741),
            data_im_out(55) => data_im_out(1773),
            data_im_out(56) => data_im_out(1805),
            data_im_out(57) => data_im_out(1837),
            data_im_out(58) => data_im_out(1869),
            data_im_out(59) => data_im_out(1901),
            data_im_out(60) => data_im_out(1933),
            data_im_out(61) => data_im_out(1965),
            data_im_out(62) => data_im_out(1997),
            data_im_out(63) => data_im_out(2029)
        );           

    URFFT_PT64_14 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(896),
            data_re_in(1) => mul_re_out(897),
            data_re_in(2) => mul_re_out(898),
            data_re_in(3) => mul_re_out(899),
            data_re_in(4) => mul_re_out(900),
            data_re_in(5) => mul_re_out(901),
            data_re_in(6) => mul_re_out(902),
            data_re_in(7) => mul_re_out(903),
            data_re_in(8) => mul_re_out(904),
            data_re_in(9) => mul_re_out(905),
            data_re_in(10) => mul_re_out(906),
            data_re_in(11) => mul_re_out(907),
            data_re_in(12) => mul_re_out(908),
            data_re_in(13) => mul_re_out(909),
            data_re_in(14) => mul_re_out(910),
            data_re_in(15) => mul_re_out(911),
            data_re_in(16) => mul_re_out(912),
            data_re_in(17) => mul_re_out(913),
            data_re_in(18) => mul_re_out(914),
            data_re_in(19) => mul_re_out(915),
            data_re_in(20) => mul_re_out(916),
            data_re_in(21) => mul_re_out(917),
            data_re_in(22) => mul_re_out(918),
            data_re_in(23) => mul_re_out(919),
            data_re_in(24) => mul_re_out(920),
            data_re_in(25) => mul_re_out(921),
            data_re_in(26) => mul_re_out(922),
            data_re_in(27) => mul_re_out(923),
            data_re_in(28) => mul_re_out(924),
            data_re_in(29) => mul_re_out(925),
            data_re_in(30) => mul_re_out(926),
            data_re_in(31) => mul_re_out(927),
            data_re_in(32) => mul_re_out(928),
            data_re_in(33) => mul_re_out(929),
            data_re_in(34) => mul_re_out(930),
            data_re_in(35) => mul_re_out(931),
            data_re_in(36) => mul_re_out(932),
            data_re_in(37) => mul_re_out(933),
            data_re_in(38) => mul_re_out(934),
            data_re_in(39) => mul_re_out(935),
            data_re_in(40) => mul_re_out(936),
            data_re_in(41) => mul_re_out(937),
            data_re_in(42) => mul_re_out(938),
            data_re_in(43) => mul_re_out(939),
            data_re_in(44) => mul_re_out(940),
            data_re_in(45) => mul_re_out(941),
            data_re_in(46) => mul_re_out(942),
            data_re_in(47) => mul_re_out(943),
            data_re_in(48) => mul_re_out(944),
            data_re_in(49) => mul_re_out(945),
            data_re_in(50) => mul_re_out(946),
            data_re_in(51) => mul_re_out(947),
            data_re_in(52) => mul_re_out(948),
            data_re_in(53) => mul_re_out(949),
            data_re_in(54) => mul_re_out(950),
            data_re_in(55) => mul_re_out(951),
            data_re_in(56) => mul_re_out(952),
            data_re_in(57) => mul_re_out(953),
            data_re_in(58) => mul_re_out(954),
            data_re_in(59) => mul_re_out(955),
            data_re_in(60) => mul_re_out(956),
            data_re_in(61) => mul_re_out(957),
            data_re_in(62) => mul_re_out(958),
            data_re_in(63) => mul_re_out(959),
            data_im_in(0) => mul_im_out(896),
            data_im_in(1) => mul_im_out(897),
            data_im_in(2) => mul_im_out(898),
            data_im_in(3) => mul_im_out(899),
            data_im_in(4) => mul_im_out(900),
            data_im_in(5) => mul_im_out(901),
            data_im_in(6) => mul_im_out(902),
            data_im_in(7) => mul_im_out(903),
            data_im_in(8) => mul_im_out(904),
            data_im_in(9) => mul_im_out(905),
            data_im_in(10) => mul_im_out(906),
            data_im_in(11) => mul_im_out(907),
            data_im_in(12) => mul_im_out(908),
            data_im_in(13) => mul_im_out(909),
            data_im_in(14) => mul_im_out(910),
            data_im_in(15) => mul_im_out(911),
            data_im_in(16) => mul_im_out(912),
            data_im_in(17) => mul_im_out(913),
            data_im_in(18) => mul_im_out(914),
            data_im_in(19) => mul_im_out(915),
            data_im_in(20) => mul_im_out(916),
            data_im_in(21) => mul_im_out(917),
            data_im_in(22) => mul_im_out(918),
            data_im_in(23) => mul_im_out(919),
            data_im_in(24) => mul_im_out(920),
            data_im_in(25) => mul_im_out(921),
            data_im_in(26) => mul_im_out(922),
            data_im_in(27) => mul_im_out(923),
            data_im_in(28) => mul_im_out(924),
            data_im_in(29) => mul_im_out(925),
            data_im_in(30) => mul_im_out(926),
            data_im_in(31) => mul_im_out(927),
            data_im_in(32) => mul_im_out(928),
            data_im_in(33) => mul_im_out(929),
            data_im_in(34) => mul_im_out(930),
            data_im_in(35) => mul_im_out(931),
            data_im_in(36) => mul_im_out(932),
            data_im_in(37) => mul_im_out(933),
            data_im_in(38) => mul_im_out(934),
            data_im_in(39) => mul_im_out(935),
            data_im_in(40) => mul_im_out(936),
            data_im_in(41) => mul_im_out(937),
            data_im_in(42) => mul_im_out(938),
            data_im_in(43) => mul_im_out(939),
            data_im_in(44) => mul_im_out(940),
            data_im_in(45) => mul_im_out(941),
            data_im_in(46) => mul_im_out(942),
            data_im_in(47) => mul_im_out(943),
            data_im_in(48) => mul_im_out(944),
            data_im_in(49) => mul_im_out(945),
            data_im_in(50) => mul_im_out(946),
            data_im_in(51) => mul_im_out(947),
            data_im_in(52) => mul_im_out(948),
            data_im_in(53) => mul_im_out(949),
            data_im_in(54) => mul_im_out(950),
            data_im_in(55) => mul_im_out(951),
            data_im_in(56) => mul_im_out(952),
            data_im_in(57) => mul_im_out(953),
            data_im_in(58) => mul_im_out(954),
            data_im_in(59) => mul_im_out(955),
            data_im_in(60) => mul_im_out(956),
            data_im_in(61) => mul_im_out(957),
            data_im_in(62) => mul_im_out(958),
            data_im_in(63) => mul_im_out(959),
            data_re_out(0) => data_re_out(14),
            data_re_out(1) => data_re_out(46),
            data_re_out(2) => data_re_out(78),
            data_re_out(3) => data_re_out(110),
            data_re_out(4) => data_re_out(142),
            data_re_out(5) => data_re_out(174),
            data_re_out(6) => data_re_out(206),
            data_re_out(7) => data_re_out(238),
            data_re_out(8) => data_re_out(270),
            data_re_out(9) => data_re_out(302),
            data_re_out(10) => data_re_out(334),
            data_re_out(11) => data_re_out(366),
            data_re_out(12) => data_re_out(398),
            data_re_out(13) => data_re_out(430),
            data_re_out(14) => data_re_out(462),
            data_re_out(15) => data_re_out(494),
            data_re_out(16) => data_re_out(526),
            data_re_out(17) => data_re_out(558),
            data_re_out(18) => data_re_out(590),
            data_re_out(19) => data_re_out(622),
            data_re_out(20) => data_re_out(654),
            data_re_out(21) => data_re_out(686),
            data_re_out(22) => data_re_out(718),
            data_re_out(23) => data_re_out(750),
            data_re_out(24) => data_re_out(782),
            data_re_out(25) => data_re_out(814),
            data_re_out(26) => data_re_out(846),
            data_re_out(27) => data_re_out(878),
            data_re_out(28) => data_re_out(910),
            data_re_out(29) => data_re_out(942),
            data_re_out(30) => data_re_out(974),
            data_re_out(31) => data_re_out(1006),
            data_re_out(32) => data_re_out(1038),
            data_re_out(33) => data_re_out(1070),
            data_re_out(34) => data_re_out(1102),
            data_re_out(35) => data_re_out(1134),
            data_re_out(36) => data_re_out(1166),
            data_re_out(37) => data_re_out(1198),
            data_re_out(38) => data_re_out(1230),
            data_re_out(39) => data_re_out(1262),
            data_re_out(40) => data_re_out(1294),
            data_re_out(41) => data_re_out(1326),
            data_re_out(42) => data_re_out(1358),
            data_re_out(43) => data_re_out(1390),
            data_re_out(44) => data_re_out(1422),
            data_re_out(45) => data_re_out(1454),
            data_re_out(46) => data_re_out(1486),
            data_re_out(47) => data_re_out(1518),
            data_re_out(48) => data_re_out(1550),
            data_re_out(49) => data_re_out(1582),
            data_re_out(50) => data_re_out(1614),
            data_re_out(51) => data_re_out(1646),
            data_re_out(52) => data_re_out(1678),
            data_re_out(53) => data_re_out(1710),
            data_re_out(54) => data_re_out(1742),
            data_re_out(55) => data_re_out(1774),
            data_re_out(56) => data_re_out(1806),
            data_re_out(57) => data_re_out(1838),
            data_re_out(58) => data_re_out(1870),
            data_re_out(59) => data_re_out(1902),
            data_re_out(60) => data_re_out(1934),
            data_re_out(61) => data_re_out(1966),
            data_re_out(62) => data_re_out(1998),
            data_re_out(63) => data_re_out(2030),
            data_im_out(0) => data_im_out(14),
            data_im_out(1) => data_im_out(46),
            data_im_out(2) => data_im_out(78),
            data_im_out(3) => data_im_out(110),
            data_im_out(4) => data_im_out(142),
            data_im_out(5) => data_im_out(174),
            data_im_out(6) => data_im_out(206),
            data_im_out(7) => data_im_out(238),
            data_im_out(8) => data_im_out(270),
            data_im_out(9) => data_im_out(302),
            data_im_out(10) => data_im_out(334),
            data_im_out(11) => data_im_out(366),
            data_im_out(12) => data_im_out(398),
            data_im_out(13) => data_im_out(430),
            data_im_out(14) => data_im_out(462),
            data_im_out(15) => data_im_out(494),
            data_im_out(16) => data_im_out(526),
            data_im_out(17) => data_im_out(558),
            data_im_out(18) => data_im_out(590),
            data_im_out(19) => data_im_out(622),
            data_im_out(20) => data_im_out(654),
            data_im_out(21) => data_im_out(686),
            data_im_out(22) => data_im_out(718),
            data_im_out(23) => data_im_out(750),
            data_im_out(24) => data_im_out(782),
            data_im_out(25) => data_im_out(814),
            data_im_out(26) => data_im_out(846),
            data_im_out(27) => data_im_out(878),
            data_im_out(28) => data_im_out(910),
            data_im_out(29) => data_im_out(942),
            data_im_out(30) => data_im_out(974),
            data_im_out(31) => data_im_out(1006),
            data_im_out(32) => data_im_out(1038),
            data_im_out(33) => data_im_out(1070),
            data_im_out(34) => data_im_out(1102),
            data_im_out(35) => data_im_out(1134),
            data_im_out(36) => data_im_out(1166),
            data_im_out(37) => data_im_out(1198),
            data_im_out(38) => data_im_out(1230),
            data_im_out(39) => data_im_out(1262),
            data_im_out(40) => data_im_out(1294),
            data_im_out(41) => data_im_out(1326),
            data_im_out(42) => data_im_out(1358),
            data_im_out(43) => data_im_out(1390),
            data_im_out(44) => data_im_out(1422),
            data_im_out(45) => data_im_out(1454),
            data_im_out(46) => data_im_out(1486),
            data_im_out(47) => data_im_out(1518),
            data_im_out(48) => data_im_out(1550),
            data_im_out(49) => data_im_out(1582),
            data_im_out(50) => data_im_out(1614),
            data_im_out(51) => data_im_out(1646),
            data_im_out(52) => data_im_out(1678),
            data_im_out(53) => data_im_out(1710),
            data_im_out(54) => data_im_out(1742),
            data_im_out(55) => data_im_out(1774),
            data_im_out(56) => data_im_out(1806),
            data_im_out(57) => data_im_out(1838),
            data_im_out(58) => data_im_out(1870),
            data_im_out(59) => data_im_out(1902),
            data_im_out(60) => data_im_out(1934),
            data_im_out(61) => data_im_out(1966),
            data_im_out(62) => data_im_out(1998),
            data_im_out(63) => data_im_out(2030)
        );           

    URFFT_PT64_15 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(960),
            data_re_in(1) => mul_re_out(961),
            data_re_in(2) => mul_re_out(962),
            data_re_in(3) => mul_re_out(963),
            data_re_in(4) => mul_re_out(964),
            data_re_in(5) => mul_re_out(965),
            data_re_in(6) => mul_re_out(966),
            data_re_in(7) => mul_re_out(967),
            data_re_in(8) => mul_re_out(968),
            data_re_in(9) => mul_re_out(969),
            data_re_in(10) => mul_re_out(970),
            data_re_in(11) => mul_re_out(971),
            data_re_in(12) => mul_re_out(972),
            data_re_in(13) => mul_re_out(973),
            data_re_in(14) => mul_re_out(974),
            data_re_in(15) => mul_re_out(975),
            data_re_in(16) => mul_re_out(976),
            data_re_in(17) => mul_re_out(977),
            data_re_in(18) => mul_re_out(978),
            data_re_in(19) => mul_re_out(979),
            data_re_in(20) => mul_re_out(980),
            data_re_in(21) => mul_re_out(981),
            data_re_in(22) => mul_re_out(982),
            data_re_in(23) => mul_re_out(983),
            data_re_in(24) => mul_re_out(984),
            data_re_in(25) => mul_re_out(985),
            data_re_in(26) => mul_re_out(986),
            data_re_in(27) => mul_re_out(987),
            data_re_in(28) => mul_re_out(988),
            data_re_in(29) => mul_re_out(989),
            data_re_in(30) => mul_re_out(990),
            data_re_in(31) => mul_re_out(991),
            data_re_in(32) => mul_re_out(992),
            data_re_in(33) => mul_re_out(993),
            data_re_in(34) => mul_re_out(994),
            data_re_in(35) => mul_re_out(995),
            data_re_in(36) => mul_re_out(996),
            data_re_in(37) => mul_re_out(997),
            data_re_in(38) => mul_re_out(998),
            data_re_in(39) => mul_re_out(999),
            data_re_in(40) => mul_re_out(1000),
            data_re_in(41) => mul_re_out(1001),
            data_re_in(42) => mul_re_out(1002),
            data_re_in(43) => mul_re_out(1003),
            data_re_in(44) => mul_re_out(1004),
            data_re_in(45) => mul_re_out(1005),
            data_re_in(46) => mul_re_out(1006),
            data_re_in(47) => mul_re_out(1007),
            data_re_in(48) => mul_re_out(1008),
            data_re_in(49) => mul_re_out(1009),
            data_re_in(50) => mul_re_out(1010),
            data_re_in(51) => mul_re_out(1011),
            data_re_in(52) => mul_re_out(1012),
            data_re_in(53) => mul_re_out(1013),
            data_re_in(54) => mul_re_out(1014),
            data_re_in(55) => mul_re_out(1015),
            data_re_in(56) => mul_re_out(1016),
            data_re_in(57) => mul_re_out(1017),
            data_re_in(58) => mul_re_out(1018),
            data_re_in(59) => mul_re_out(1019),
            data_re_in(60) => mul_re_out(1020),
            data_re_in(61) => mul_re_out(1021),
            data_re_in(62) => mul_re_out(1022),
            data_re_in(63) => mul_re_out(1023),
            data_im_in(0) => mul_im_out(960),
            data_im_in(1) => mul_im_out(961),
            data_im_in(2) => mul_im_out(962),
            data_im_in(3) => mul_im_out(963),
            data_im_in(4) => mul_im_out(964),
            data_im_in(5) => mul_im_out(965),
            data_im_in(6) => mul_im_out(966),
            data_im_in(7) => mul_im_out(967),
            data_im_in(8) => mul_im_out(968),
            data_im_in(9) => mul_im_out(969),
            data_im_in(10) => mul_im_out(970),
            data_im_in(11) => mul_im_out(971),
            data_im_in(12) => mul_im_out(972),
            data_im_in(13) => mul_im_out(973),
            data_im_in(14) => mul_im_out(974),
            data_im_in(15) => mul_im_out(975),
            data_im_in(16) => mul_im_out(976),
            data_im_in(17) => mul_im_out(977),
            data_im_in(18) => mul_im_out(978),
            data_im_in(19) => mul_im_out(979),
            data_im_in(20) => mul_im_out(980),
            data_im_in(21) => mul_im_out(981),
            data_im_in(22) => mul_im_out(982),
            data_im_in(23) => mul_im_out(983),
            data_im_in(24) => mul_im_out(984),
            data_im_in(25) => mul_im_out(985),
            data_im_in(26) => mul_im_out(986),
            data_im_in(27) => mul_im_out(987),
            data_im_in(28) => mul_im_out(988),
            data_im_in(29) => mul_im_out(989),
            data_im_in(30) => mul_im_out(990),
            data_im_in(31) => mul_im_out(991),
            data_im_in(32) => mul_im_out(992),
            data_im_in(33) => mul_im_out(993),
            data_im_in(34) => mul_im_out(994),
            data_im_in(35) => mul_im_out(995),
            data_im_in(36) => mul_im_out(996),
            data_im_in(37) => mul_im_out(997),
            data_im_in(38) => mul_im_out(998),
            data_im_in(39) => mul_im_out(999),
            data_im_in(40) => mul_im_out(1000),
            data_im_in(41) => mul_im_out(1001),
            data_im_in(42) => mul_im_out(1002),
            data_im_in(43) => mul_im_out(1003),
            data_im_in(44) => mul_im_out(1004),
            data_im_in(45) => mul_im_out(1005),
            data_im_in(46) => mul_im_out(1006),
            data_im_in(47) => mul_im_out(1007),
            data_im_in(48) => mul_im_out(1008),
            data_im_in(49) => mul_im_out(1009),
            data_im_in(50) => mul_im_out(1010),
            data_im_in(51) => mul_im_out(1011),
            data_im_in(52) => mul_im_out(1012),
            data_im_in(53) => mul_im_out(1013),
            data_im_in(54) => mul_im_out(1014),
            data_im_in(55) => mul_im_out(1015),
            data_im_in(56) => mul_im_out(1016),
            data_im_in(57) => mul_im_out(1017),
            data_im_in(58) => mul_im_out(1018),
            data_im_in(59) => mul_im_out(1019),
            data_im_in(60) => mul_im_out(1020),
            data_im_in(61) => mul_im_out(1021),
            data_im_in(62) => mul_im_out(1022),
            data_im_in(63) => mul_im_out(1023),
            data_re_out(0) => data_re_out(15),
            data_re_out(1) => data_re_out(47),
            data_re_out(2) => data_re_out(79),
            data_re_out(3) => data_re_out(111),
            data_re_out(4) => data_re_out(143),
            data_re_out(5) => data_re_out(175),
            data_re_out(6) => data_re_out(207),
            data_re_out(7) => data_re_out(239),
            data_re_out(8) => data_re_out(271),
            data_re_out(9) => data_re_out(303),
            data_re_out(10) => data_re_out(335),
            data_re_out(11) => data_re_out(367),
            data_re_out(12) => data_re_out(399),
            data_re_out(13) => data_re_out(431),
            data_re_out(14) => data_re_out(463),
            data_re_out(15) => data_re_out(495),
            data_re_out(16) => data_re_out(527),
            data_re_out(17) => data_re_out(559),
            data_re_out(18) => data_re_out(591),
            data_re_out(19) => data_re_out(623),
            data_re_out(20) => data_re_out(655),
            data_re_out(21) => data_re_out(687),
            data_re_out(22) => data_re_out(719),
            data_re_out(23) => data_re_out(751),
            data_re_out(24) => data_re_out(783),
            data_re_out(25) => data_re_out(815),
            data_re_out(26) => data_re_out(847),
            data_re_out(27) => data_re_out(879),
            data_re_out(28) => data_re_out(911),
            data_re_out(29) => data_re_out(943),
            data_re_out(30) => data_re_out(975),
            data_re_out(31) => data_re_out(1007),
            data_re_out(32) => data_re_out(1039),
            data_re_out(33) => data_re_out(1071),
            data_re_out(34) => data_re_out(1103),
            data_re_out(35) => data_re_out(1135),
            data_re_out(36) => data_re_out(1167),
            data_re_out(37) => data_re_out(1199),
            data_re_out(38) => data_re_out(1231),
            data_re_out(39) => data_re_out(1263),
            data_re_out(40) => data_re_out(1295),
            data_re_out(41) => data_re_out(1327),
            data_re_out(42) => data_re_out(1359),
            data_re_out(43) => data_re_out(1391),
            data_re_out(44) => data_re_out(1423),
            data_re_out(45) => data_re_out(1455),
            data_re_out(46) => data_re_out(1487),
            data_re_out(47) => data_re_out(1519),
            data_re_out(48) => data_re_out(1551),
            data_re_out(49) => data_re_out(1583),
            data_re_out(50) => data_re_out(1615),
            data_re_out(51) => data_re_out(1647),
            data_re_out(52) => data_re_out(1679),
            data_re_out(53) => data_re_out(1711),
            data_re_out(54) => data_re_out(1743),
            data_re_out(55) => data_re_out(1775),
            data_re_out(56) => data_re_out(1807),
            data_re_out(57) => data_re_out(1839),
            data_re_out(58) => data_re_out(1871),
            data_re_out(59) => data_re_out(1903),
            data_re_out(60) => data_re_out(1935),
            data_re_out(61) => data_re_out(1967),
            data_re_out(62) => data_re_out(1999),
            data_re_out(63) => data_re_out(2031),
            data_im_out(0) => data_im_out(15),
            data_im_out(1) => data_im_out(47),
            data_im_out(2) => data_im_out(79),
            data_im_out(3) => data_im_out(111),
            data_im_out(4) => data_im_out(143),
            data_im_out(5) => data_im_out(175),
            data_im_out(6) => data_im_out(207),
            data_im_out(7) => data_im_out(239),
            data_im_out(8) => data_im_out(271),
            data_im_out(9) => data_im_out(303),
            data_im_out(10) => data_im_out(335),
            data_im_out(11) => data_im_out(367),
            data_im_out(12) => data_im_out(399),
            data_im_out(13) => data_im_out(431),
            data_im_out(14) => data_im_out(463),
            data_im_out(15) => data_im_out(495),
            data_im_out(16) => data_im_out(527),
            data_im_out(17) => data_im_out(559),
            data_im_out(18) => data_im_out(591),
            data_im_out(19) => data_im_out(623),
            data_im_out(20) => data_im_out(655),
            data_im_out(21) => data_im_out(687),
            data_im_out(22) => data_im_out(719),
            data_im_out(23) => data_im_out(751),
            data_im_out(24) => data_im_out(783),
            data_im_out(25) => data_im_out(815),
            data_im_out(26) => data_im_out(847),
            data_im_out(27) => data_im_out(879),
            data_im_out(28) => data_im_out(911),
            data_im_out(29) => data_im_out(943),
            data_im_out(30) => data_im_out(975),
            data_im_out(31) => data_im_out(1007),
            data_im_out(32) => data_im_out(1039),
            data_im_out(33) => data_im_out(1071),
            data_im_out(34) => data_im_out(1103),
            data_im_out(35) => data_im_out(1135),
            data_im_out(36) => data_im_out(1167),
            data_im_out(37) => data_im_out(1199),
            data_im_out(38) => data_im_out(1231),
            data_im_out(39) => data_im_out(1263),
            data_im_out(40) => data_im_out(1295),
            data_im_out(41) => data_im_out(1327),
            data_im_out(42) => data_im_out(1359),
            data_im_out(43) => data_im_out(1391),
            data_im_out(44) => data_im_out(1423),
            data_im_out(45) => data_im_out(1455),
            data_im_out(46) => data_im_out(1487),
            data_im_out(47) => data_im_out(1519),
            data_im_out(48) => data_im_out(1551),
            data_im_out(49) => data_im_out(1583),
            data_im_out(50) => data_im_out(1615),
            data_im_out(51) => data_im_out(1647),
            data_im_out(52) => data_im_out(1679),
            data_im_out(53) => data_im_out(1711),
            data_im_out(54) => data_im_out(1743),
            data_im_out(55) => data_im_out(1775),
            data_im_out(56) => data_im_out(1807),
            data_im_out(57) => data_im_out(1839),
            data_im_out(58) => data_im_out(1871),
            data_im_out(59) => data_im_out(1903),
            data_im_out(60) => data_im_out(1935),
            data_im_out(61) => data_im_out(1967),
            data_im_out(62) => data_im_out(1999),
            data_im_out(63) => data_im_out(2031)
        );           

    URFFT_PT64_16 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1024),
            data_re_in(1) => mul_re_out(1025),
            data_re_in(2) => mul_re_out(1026),
            data_re_in(3) => mul_re_out(1027),
            data_re_in(4) => mul_re_out(1028),
            data_re_in(5) => mul_re_out(1029),
            data_re_in(6) => mul_re_out(1030),
            data_re_in(7) => mul_re_out(1031),
            data_re_in(8) => mul_re_out(1032),
            data_re_in(9) => mul_re_out(1033),
            data_re_in(10) => mul_re_out(1034),
            data_re_in(11) => mul_re_out(1035),
            data_re_in(12) => mul_re_out(1036),
            data_re_in(13) => mul_re_out(1037),
            data_re_in(14) => mul_re_out(1038),
            data_re_in(15) => mul_re_out(1039),
            data_re_in(16) => mul_re_out(1040),
            data_re_in(17) => mul_re_out(1041),
            data_re_in(18) => mul_re_out(1042),
            data_re_in(19) => mul_re_out(1043),
            data_re_in(20) => mul_re_out(1044),
            data_re_in(21) => mul_re_out(1045),
            data_re_in(22) => mul_re_out(1046),
            data_re_in(23) => mul_re_out(1047),
            data_re_in(24) => mul_re_out(1048),
            data_re_in(25) => mul_re_out(1049),
            data_re_in(26) => mul_re_out(1050),
            data_re_in(27) => mul_re_out(1051),
            data_re_in(28) => mul_re_out(1052),
            data_re_in(29) => mul_re_out(1053),
            data_re_in(30) => mul_re_out(1054),
            data_re_in(31) => mul_re_out(1055),
            data_re_in(32) => mul_re_out(1056),
            data_re_in(33) => mul_re_out(1057),
            data_re_in(34) => mul_re_out(1058),
            data_re_in(35) => mul_re_out(1059),
            data_re_in(36) => mul_re_out(1060),
            data_re_in(37) => mul_re_out(1061),
            data_re_in(38) => mul_re_out(1062),
            data_re_in(39) => mul_re_out(1063),
            data_re_in(40) => mul_re_out(1064),
            data_re_in(41) => mul_re_out(1065),
            data_re_in(42) => mul_re_out(1066),
            data_re_in(43) => mul_re_out(1067),
            data_re_in(44) => mul_re_out(1068),
            data_re_in(45) => mul_re_out(1069),
            data_re_in(46) => mul_re_out(1070),
            data_re_in(47) => mul_re_out(1071),
            data_re_in(48) => mul_re_out(1072),
            data_re_in(49) => mul_re_out(1073),
            data_re_in(50) => mul_re_out(1074),
            data_re_in(51) => mul_re_out(1075),
            data_re_in(52) => mul_re_out(1076),
            data_re_in(53) => mul_re_out(1077),
            data_re_in(54) => mul_re_out(1078),
            data_re_in(55) => mul_re_out(1079),
            data_re_in(56) => mul_re_out(1080),
            data_re_in(57) => mul_re_out(1081),
            data_re_in(58) => mul_re_out(1082),
            data_re_in(59) => mul_re_out(1083),
            data_re_in(60) => mul_re_out(1084),
            data_re_in(61) => mul_re_out(1085),
            data_re_in(62) => mul_re_out(1086),
            data_re_in(63) => mul_re_out(1087),
            data_im_in(0) => mul_im_out(1024),
            data_im_in(1) => mul_im_out(1025),
            data_im_in(2) => mul_im_out(1026),
            data_im_in(3) => mul_im_out(1027),
            data_im_in(4) => mul_im_out(1028),
            data_im_in(5) => mul_im_out(1029),
            data_im_in(6) => mul_im_out(1030),
            data_im_in(7) => mul_im_out(1031),
            data_im_in(8) => mul_im_out(1032),
            data_im_in(9) => mul_im_out(1033),
            data_im_in(10) => mul_im_out(1034),
            data_im_in(11) => mul_im_out(1035),
            data_im_in(12) => mul_im_out(1036),
            data_im_in(13) => mul_im_out(1037),
            data_im_in(14) => mul_im_out(1038),
            data_im_in(15) => mul_im_out(1039),
            data_im_in(16) => mul_im_out(1040),
            data_im_in(17) => mul_im_out(1041),
            data_im_in(18) => mul_im_out(1042),
            data_im_in(19) => mul_im_out(1043),
            data_im_in(20) => mul_im_out(1044),
            data_im_in(21) => mul_im_out(1045),
            data_im_in(22) => mul_im_out(1046),
            data_im_in(23) => mul_im_out(1047),
            data_im_in(24) => mul_im_out(1048),
            data_im_in(25) => mul_im_out(1049),
            data_im_in(26) => mul_im_out(1050),
            data_im_in(27) => mul_im_out(1051),
            data_im_in(28) => mul_im_out(1052),
            data_im_in(29) => mul_im_out(1053),
            data_im_in(30) => mul_im_out(1054),
            data_im_in(31) => mul_im_out(1055),
            data_im_in(32) => mul_im_out(1056),
            data_im_in(33) => mul_im_out(1057),
            data_im_in(34) => mul_im_out(1058),
            data_im_in(35) => mul_im_out(1059),
            data_im_in(36) => mul_im_out(1060),
            data_im_in(37) => mul_im_out(1061),
            data_im_in(38) => mul_im_out(1062),
            data_im_in(39) => mul_im_out(1063),
            data_im_in(40) => mul_im_out(1064),
            data_im_in(41) => mul_im_out(1065),
            data_im_in(42) => mul_im_out(1066),
            data_im_in(43) => mul_im_out(1067),
            data_im_in(44) => mul_im_out(1068),
            data_im_in(45) => mul_im_out(1069),
            data_im_in(46) => mul_im_out(1070),
            data_im_in(47) => mul_im_out(1071),
            data_im_in(48) => mul_im_out(1072),
            data_im_in(49) => mul_im_out(1073),
            data_im_in(50) => mul_im_out(1074),
            data_im_in(51) => mul_im_out(1075),
            data_im_in(52) => mul_im_out(1076),
            data_im_in(53) => mul_im_out(1077),
            data_im_in(54) => mul_im_out(1078),
            data_im_in(55) => mul_im_out(1079),
            data_im_in(56) => mul_im_out(1080),
            data_im_in(57) => mul_im_out(1081),
            data_im_in(58) => mul_im_out(1082),
            data_im_in(59) => mul_im_out(1083),
            data_im_in(60) => mul_im_out(1084),
            data_im_in(61) => mul_im_out(1085),
            data_im_in(62) => mul_im_out(1086),
            data_im_in(63) => mul_im_out(1087),
            data_re_out(0) => data_re_out(16),
            data_re_out(1) => data_re_out(48),
            data_re_out(2) => data_re_out(80),
            data_re_out(3) => data_re_out(112),
            data_re_out(4) => data_re_out(144),
            data_re_out(5) => data_re_out(176),
            data_re_out(6) => data_re_out(208),
            data_re_out(7) => data_re_out(240),
            data_re_out(8) => data_re_out(272),
            data_re_out(9) => data_re_out(304),
            data_re_out(10) => data_re_out(336),
            data_re_out(11) => data_re_out(368),
            data_re_out(12) => data_re_out(400),
            data_re_out(13) => data_re_out(432),
            data_re_out(14) => data_re_out(464),
            data_re_out(15) => data_re_out(496),
            data_re_out(16) => data_re_out(528),
            data_re_out(17) => data_re_out(560),
            data_re_out(18) => data_re_out(592),
            data_re_out(19) => data_re_out(624),
            data_re_out(20) => data_re_out(656),
            data_re_out(21) => data_re_out(688),
            data_re_out(22) => data_re_out(720),
            data_re_out(23) => data_re_out(752),
            data_re_out(24) => data_re_out(784),
            data_re_out(25) => data_re_out(816),
            data_re_out(26) => data_re_out(848),
            data_re_out(27) => data_re_out(880),
            data_re_out(28) => data_re_out(912),
            data_re_out(29) => data_re_out(944),
            data_re_out(30) => data_re_out(976),
            data_re_out(31) => data_re_out(1008),
            data_re_out(32) => data_re_out(1040),
            data_re_out(33) => data_re_out(1072),
            data_re_out(34) => data_re_out(1104),
            data_re_out(35) => data_re_out(1136),
            data_re_out(36) => data_re_out(1168),
            data_re_out(37) => data_re_out(1200),
            data_re_out(38) => data_re_out(1232),
            data_re_out(39) => data_re_out(1264),
            data_re_out(40) => data_re_out(1296),
            data_re_out(41) => data_re_out(1328),
            data_re_out(42) => data_re_out(1360),
            data_re_out(43) => data_re_out(1392),
            data_re_out(44) => data_re_out(1424),
            data_re_out(45) => data_re_out(1456),
            data_re_out(46) => data_re_out(1488),
            data_re_out(47) => data_re_out(1520),
            data_re_out(48) => data_re_out(1552),
            data_re_out(49) => data_re_out(1584),
            data_re_out(50) => data_re_out(1616),
            data_re_out(51) => data_re_out(1648),
            data_re_out(52) => data_re_out(1680),
            data_re_out(53) => data_re_out(1712),
            data_re_out(54) => data_re_out(1744),
            data_re_out(55) => data_re_out(1776),
            data_re_out(56) => data_re_out(1808),
            data_re_out(57) => data_re_out(1840),
            data_re_out(58) => data_re_out(1872),
            data_re_out(59) => data_re_out(1904),
            data_re_out(60) => data_re_out(1936),
            data_re_out(61) => data_re_out(1968),
            data_re_out(62) => data_re_out(2000),
            data_re_out(63) => data_re_out(2032),
            data_im_out(0) => data_im_out(16),
            data_im_out(1) => data_im_out(48),
            data_im_out(2) => data_im_out(80),
            data_im_out(3) => data_im_out(112),
            data_im_out(4) => data_im_out(144),
            data_im_out(5) => data_im_out(176),
            data_im_out(6) => data_im_out(208),
            data_im_out(7) => data_im_out(240),
            data_im_out(8) => data_im_out(272),
            data_im_out(9) => data_im_out(304),
            data_im_out(10) => data_im_out(336),
            data_im_out(11) => data_im_out(368),
            data_im_out(12) => data_im_out(400),
            data_im_out(13) => data_im_out(432),
            data_im_out(14) => data_im_out(464),
            data_im_out(15) => data_im_out(496),
            data_im_out(16) => data_im_out(528),
            data_im_out(17) => data_im_out(560),
            data_im_out(18) => data_im_out(592),
            data_im_out(19) => data_im_out(624),
            data_im_out(20) => data_im_out(656),
            data_im_out(21) => data_im_out(688),
            data_im_out(22) => data_im_out(720),
            data_im_out(23) => data_im_out(752),
            data_im_out(24) => data_im_out(784),
            data_im_out(25) => data_im_out(816),
            data_im_out(26) => data_im_out(848),
            data_im_out(27) => data_im_out(880),
            data_im_out(28) => data_im_out(912),
            data_im_out(29) => data_im_out(944),
            data_im_out(30) => data_im_out(976),
            data_im_out(31) => data_im_out(1008),
            data_im_out(32) => data_im_out(1040),
            data_im_out(33) => data_im_out(1072),
            data_im_out(34) => data_im_out(1104),
            data_im_out(35) => data_im_out(1136),
            data_im_out(36) => data_im_out(1168),
            data_im_out(37) => data_im_out(1200),
            data_im_out(38) => data_im_out(1232),
            data_im_out(39) => data_im_out(1264),
            data_im_out(40) => data_im_out(1296),
            data_im_out(41) => data_im_out(1328),
            data_im_out(42) => data_im_out(1360),
            data_im_out(43) => data_im_out(1392),
            data_im_out(44) => data_im_out(1424),
            data_im_out(45) => data_im_out(1456),
            data_im_out(46) => data_im_out(1488),
            data_im_out(47) => data_im_out(1520),
            data_im_out(48) => data_im_out(1552),
            data_im_out(49) => data_im_out(1584),
            data_im_out(50) => data_im_out(1616),
            data_im_out(51) => data_im_out(1648),
            data_im_out(52) => data_im_out(1680),
            data_im_out(53) => data_im_out(1712),
            data_im_out(54) => data_im_out(1744),
            data_im_out(55) => data_im_out(1776),
            data_im_out(56) => data_im_out(1808),
            data_im_out(57) => data_im_out(1840),
            data_im_out(58) => data_im_out(1872),
            data_im_out(59) => data_im_out(1904),
            data_im_out(60) => data_im_out(1936),
            data_im_out(61) => data_im_out(1968),
            data_im_out(62) => data_im_out(2000),
            data_im_out(63) => data_im_out(2032)
        );           

    URFFT_PT64_17 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1088),
            data_re_in(1) => mul_re_out(1089),
            data_re_in(2) => mul_re_out(1090),
            data_re_in(3) => mul_re_out(1091),
            data_re_in(4) => mul_re_out(1092),
            data_re_in(5) => mul_re_out(1093),
            data_re_in(6) => mul_re_out(1094),
            data_re_in(7) => mul_re_out(1095),
            data_re_in(8) => mul_re_out(1096),
            data_re_in(9) => mul_re_out(1097),
            data_re_in(10) => mul_re_out(1098),
            data_re_in(11) => mul_re_out(1099),
            data_re_in(12) => mul_re_out(1100),
            data_re_in(13) => mul_re_out(1101),
            data_re_in(14) => mul_re_out(1102),
            data_re_in(15) => mul_re_out(1103),
            data_re_in(16) => mul_re_out(1104),
            data_re_in(17) => mul_re_out(1105),
            data_re_in(18) => mul_re_out(1106),
            data_re_in(19) => mul_re_out(1107),
            data_re_in(20) => mul_re_out(1108),
            data_re_in(21) => mul_re_out(1109),
            data_re_in(22) => mul_re_out(1110),
            data_re_in(23) => mul_re_out(1111),
            data_re_in(24) => mul_re_out(1112),
            data_re_in(25) => mul_re_out(1113),
            data_re_in(26) => mul_re_out(1114),
            data_re_in(27) => mul_re_out(1115),
            data_re_in(28) => mul_re_out(1116),
            data_re_in(29) => mul_re_out(1117),
            data_re_in(30) => mul_re_out(1118),
            data_re_in(31) => mul_re_out(1119),
            data_re_in(32) => mul_re_out(1120),
            data_re_in(33) => mul_re_out(1121),
            data_re_in(34) => mul_re_out(1122),
            data_re_in(35) => mul_re_out(1123),
            data_re_in(36) => mul_re_out(1124),
            data_re_in(37) => mul_re_out(1125),
            data_re_in(38) => mul_re_out(1126),
            data_re_in(39) => mul_re_out(1127),
            data_re_in(40) => mul_re_out(1128),
            data_re_in(41) => mul_re_out(1129),
            data_re_in(42) => mul_re_out(1130),
            data_re_in(43) => mul_re_out(1131),
            data_re_in(44) => mul_re_out(1132),
            data_re_in(45) => mul_re_out(1133),
            data_re_in(46) => mul_re_out(1134),
            data_re_in(47) => mul_re_out(1135),
            data_re_in(48) => mul_re_out(1136),
            data_re_in(49) => mul_re_out(1137),
            data_re_in(50) => mul_re_out(1138),
            data_re_in(51) => mul_re_out(1139),
            data_re_in(52) => mul_re_out(1140),
            data_re_in(53) => mul_re_out(1141),
            data_re_in(54) => mul_re_out(1142),
            data_re_in(55) => mul_re_out(1143),
            data_re_in(56) => mul_re_out(1144),
            data_re_in(57) => mul_re_out(1145),
            data_re_in(58) => mul_re_out(1146),
            data_re_in(59) => mul_re_out(1147),
            data_re_in(60) => mul_re_out(1148),
            data_re_in(61) => mul_re_out(1149),
            data_re_in(62) => mul_re_out(1150),
            data_re_in(63) => mul_re_out(1151),
            data_im_in(0) => mul_im_out(1088),
            data_im_in(1) => mul_im_out(1089),
            data_im_in(2) => mul_im_out(1090),
            data_im_in(3) => mul_im_out(1091),
            data_im_in(4) => mul_im_out(1092),
            data_im_in(5) => mul_im_out(1093),
            data_im_in(6) => mul_im_out(1094),
            data_im_in(7) => mul_im_out(1095),
            data_im_in(8) => mul_im_out(1096),
            data_im_in(9) => mul_im_out(1097),
            data_im_in(10) => mul_im_out(1098),
            data_im_in(11) => mul_im_out(1099),
            data_im_in(12) => mul_im_out(1100),
            data_im_in(13) => mul_im_out(1101),
            data_im_in(14) => mul_im_out(1102),
            data_im_in(15) => mul_im_out(1103),
            data_im_in(16) => mul_im_out(1104),
            data_im_in(17) => mul_im_out(1105),
            data_im_in(18) => mul_im_out(1106),
            data_im_in(19) => mul_im_out(1107),
            data_im_in(20) => mul_im_out(1108),
            data_im_in(21) => mul_im_out(1109),
            data_im_in(22) => mul_im_out(1110),
            data_im_in(23) => mul_im_out(1111),
            data_im_in(24) => mul_im_out(1112),
            data_im_in(25) => mul_im_out(1113),
            data_im_in(26) => mul_im_out(1114),
            data_im_in(27) => mul_im_out(1115),
            data_im_in(28) => mul_im_out(1116),
            data_im_in(29) => mul_im_out(1117),
            data_im_in(30) => mul_im_out(1118),
            data_im_in(31) => mul_im_out(1119),
            data_im_in(32) => mul_im_out(1120),
            data_im_in(33) => mul_im_out(1121),
            data_im_in(34) => mul_im_out(1122),
            data_im_in(35) => mul_im_out(1123),
            data_im_in(36) => mul_im_out(1124),
            data_im_in(37) => mul_im_out(1125),
            data_im_in(38) => mul_im_out(1126),
            data_im_in(39) => mul_im_out(1127),
            data_im_in(40) => mul_im_out(1128),
            data_im_in(41) => mul_im_out(1129),
            data_im_in(42) => mul_im_out(1130),
            data_im_in(43) => mul_im_out(1131),
            data_im_in(44) => mul_im_out(1132),
            data_im_in(45) => mul_im_out(1133),
            data_im_in(46) => mul_im_out(1134),
            data_im_in(47) => mul_im_out(1135),
            data_im_in(48) => mul_im_out(1136),
            data_im_in(49) => mul_im_out(1137),
            data_im_in(50) => mul_im_out(1138),
            data_im_in(51) => mul_im_out(1139),
            data_im_in(52) => mul_im_out(1140),
            data_im_in(53) => mul_im_out(1141),
            data_im_in(54) => mul_im_out(1142),
            data_im_in(55) => mul_im_out(1143),
            data_im_in(56) => mul_im_out(1144),
            data_im_in(57) => mul_im_out(1145),
            data_im_in(58) => mul_im_out(1146),
            data_im_in(59) => mul_im_out(1147),
            data_im_in(60) => mul_im_out(1148),
            data_im_in(61) => mul_im_out(1149),
            data_im_in(62) => mul_im_out(1150),
            data_im_in(63) => mul_im_out(1151),
            data_re_out(0) => data_re_out(17),
            data_re_out(1) => data_re_out(49),
            data_re_out(2) => data_re_out(81),
            data_re_out(3) => data_re_out(113),
            data_re_out(4) => data_re_out(145),
            data_re_out(5) => data_re_out(177),
            data_re_out(6) => data_re_out(209),
            data_re_out(7) => data_re_out(241),
            data_re_out(8) => data_re_out(273),
            data_re_out(9) => data_re_out(305),
            data_re_out(10) => data_re_out(337),
            data_re_out(11) => data_re_out(369),
            data_re_out(12) => data_re_out(401),
            data_re_out(13) => data_re_out(433),
            data_re_out(14) => data_re_out(465),
            data_re_out(15) => data_re_out(497),
            data_re_out(16) => data_re_out(529),
            data_re_out(17) => data_re_out(561),
            data_re_out(18) => data_re_out(593),
            data_re_out(19) => data_re_out(625),
            data_re_out(20) => data_re_out(657),
            data_re_out(21) => data_re_out(689),
            data_re_out(22) => data_re_out(721),
            data_re_out(23) => data_re_out(753),
            data_re_out(24) => data_re_out(785),
            data_re_out(25) => data_re_out(817),
            data_re_out(26) => data_re_out(849),
            data_re_out(27) => data_re_out(881),
            data_re_out(28) => data_re_out(913),
            data_re_out(29) => data_re_out(945),
            data_re_out(30) => data_re_out(977),
            data_re_out(31) => data_re_out(1009),
            data_re_out(32) => data_re_out(1041),
            data_re_out(33) => data_re_out(1073),
            data_re_out(34) => data_re_out(1105),
            data_re_out(35) => data_re_out(1137),
            data_re_out(36) => data_re_out(1169),
            data_re_out(37) => data_re_out(1201),
            data_re_out(38) => data_re_out(1233),
            data_re_out(39) => data_re_out(1265),
            data_re_out(40) => data_re_out(1297),
            data_re_out(41) => data_re_out(1329),
            data_re_out(42) => data_re_out(1361),
            data_re_out(43) => data_re_out(1393),
            data_re_out(44) => data_re_out(1425),
            data_re_out(45) => data_re_out(1457),
            data_re_out(46) => data_re_out(1489),
            data_re_out(47) => data_re_out(1521),
            data_re_out(48) => data_re_out(1553),
            data_re_out(49) => data_re_out(1585),
            data_re_out(50) => data_re_out(1617),
            data_re_out(51) => data_re_out(1649),
            data_re_out(52) => data_re_out(1681),
            data_re_out(53) => data_re_out(1713),
            data_re_out(54) => data_re_out(1745),
            data_re_out(55) => data_re_out(1777),
            data_re_out(56) => data_re_out(1809),
            data_re_out(57) => data_re_out(1841),
            data_re_out(58) => data_re_out(1873),
            data_re_out(59) => data_re_out(1905),
            data_re_out(60) => data_re_out(1937),
            data_re_out(61) => data_re_out(1969),
            data_re_out(62) => data_re_out(2001),
            data_re_out(63) => data_re_out(2033),
            data_im_out(0) => data_im_out(17),
            data_im_out(1) => data_im_out(49),
            data_im_out(2) => data_im_out(81),
            data_im_out(3) => data_im_out(113),
            data_im_out(4) => data_im_out(145),
            data_im_out(5) => data_im_out(177),
            data_im_out(6) => data_im_out(209),
            data_im_out(7) => data_im_out(241),
            data_im_out(8) => data_im_out(273),
            data_im_out(9) => data_im_out(305),
            data_im_out(10) => data_im_out(337),
            data_im_out(11) => data_im_out(369),
            data_im_out(12) => data_im_out(401),
            data_im_out(13) => data_im_out(433),
            data_im_out(14) => data_im_out(465),
            data_im_out(15) => data_im_out(497),
            data_im_out(16) => data_im_out(529),
            data_im_out(17) => data_im_out(561),
            data_im_out(18) => data_im_out(593),
            data_im_out(19) => data_im_out(625),
            data_im_out(20) => data_im_out(657),
            data_im_out(21) => data_im_out(689),
            data_im_out(22) => data_im_out(721),
            data_im_out(23) => data_im_out(753),
            data_im_out(24) => data_im_out(785),
            data_im_out(25) => data_im_out(817),
            data_im_out(26) => data_im_out(849),
            data_im_out(27) => data_im_out(881),
            data_im_out(28) => data_im_out(913),
            data_im_out(29) => data_im_out(945),
            data_im_out(30) => data_im_out(977),
            data_im_out(31) => data_im_out(1009),
            data_im_out(32) => data_im_out(1041),
            data_im_out(33) => data_im_out(1073),
            data_im_out(34) => data_im_out(1105),
            data_im_out(35) => data_im_out(1137),
            data_im_out(36) => data_im_out(1169),
            data_im_out(37) => data_im_out(1201),
            data_im_out(38) => data_im_out(1233),
            data_im_out(39) => data_im_out(1265),
            data_im_out(40) => data_im_out(1297),
            data_im_out(41) => data_im_out(1329),
            data_im_out(42) => data_im_out(1361),
            data_im_out(43) => data_im_out(1393),
            data_im_out(44) => data_im_out(1425),
            data_im_out(45) => data_im_out(1457),
            data_im_out(46) => data_im_out(1489),
            data_im_out(47) => data_im_out(1521),
            data_im_out(48) => data_im_out(1553),
            data_im_out(49) => data_im_out(1585),
            data_im_out(50) => data_im_out(1617),
            data_im_out(51) => data_im_out(1649),
            data_im_out(52) => data_im_out(1681),
            data_im_out(53) => data_im_out(1713),
            data_im_out(54) => data_im_out(1745),
            data_im_out(55) => data_im_out(1777),
            data_im_out(56) => data_im_out(1809),
            data_im_out(57) => data_im_out(1841),
            data_im_out(58) => data_im_out(1873),
            data_im_out(59) => data_im_out(1905),
            data_im_out(60) => data_im_out(1937),
            data_im_out(61) => data_im_out(1969),
            data_im_out(62) => data_im_out(2001),
            data_im_out(63) => data_im_out(2033)
        );           

    URFFT_PT64_18 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1152),
            data_re_in(1) => mul_re_out(1153),
            data_re_in(2) => mul_re_out(1154),
            data_re_in(3) => mul_re_out(1155),
            data_re_in(4) => mul_re_out(1156),
            data_re_in(5) => mul_re_out(1157),
            data_re_in(6) => mul_re_out(1158),
            data_re_in(7) => mul_re_out(1159),
            data_re_in(8) => mul_re_out(1160),
            data_re_in(9) => mul_re_out(1161),
            data_re_in(10) => mul_re_out(1162),
            data_re_in(11) => mul_re_out(1163),
            data_re_in(12) => mul_re_out(1164),
            data_re_in(13) => mul_re_out(1165),
            data_re_in(14) => mul_re_out(1166),
            data_re_in(15) => mul_re_out(1167),
            data_re_in(16) => mul_re_out(1168),
            data_re_in(17) => mul_re_out(1169),
            data_re_in(18) => mul_re_out(1170),
            data_re_in(19) => mul_re_out(1171),
            data_re_in(20) => mul_re_out(1172),
            data_re_in(21) => mul_re_out(1173),
            data_re_in(22) => mul_re_out(1174),
            data_re_in(23) => mul_re_out(1175),
            data_re_in(24) => mul_re_out(1176),
            data_re_in(25) => mul_re_out(1177),
            data_re_in(26) => mul_re_out(1178),
            data_re_in(27) => mul_re_out(1179),
            data_re_in(28) => mul_re_out(1180),
            data_re_in(29) => mul_re_out(1181),
            data_re_in(30) => mul_re_out(1182),
            data_re_in(31) => mul_re_out(1183),
            data_re_in(32) => mul_re_out(1184),
            data_re_in(33) => mul_re_out(1185),
            data_re_in(34) => mul_re_out(1186),
            data_re_in(35) => mul_re_out(1187),
            data_re_in(36) => mul_re_out(1188),
            data_re_in(37) => mul_re_out(1189),
            data_re_in(38) => mul_re_out(1190),
            data_re_in(39) => mul_re_out(1191),
            data_re_in(40) => mul_re_out(1192),
            data_re_in(41) => mul_re_out(1193),
            data_re_in(42) => mul_re_out(1194),
            data_re_in(43) => mul_re_out(1195),
            data_re_in(44) => mul_re_out(1196),
            data_re_in(45) => mul_re_out(1197),
            data_re_in(46) => mul_re_out(1198),
            data_re_in(47) => mul_re_out(1199),
            data_re_in(48) => mul_re_out(1200),
            data_re_in(49) => mul_re_out(1201),
            data_re_in(50) => mul_re_out(1202),
            data_re_in(51) => mul_re_out(1203),
            data_re_in(52) => mul_re_out(1204),
            data_re_in(53) => mul_re_out(1205),
            data_re_in(54) => mul_re_out(1206),
            data_re_in(55) => mul_re_out(1207),
            data_re_in(56) => mul_re_out(1208),
            data_re_in(57) => mul_re_out(1209),
            data_re_in(58) => mul_re_out(1210),
            data_re_in(59) => mul_re_out(1211),
            data_re_in(60) => mul_re_out(1212),
            data_re_in(61) => mul_re_out(1213),
            data_re_in(62) => mul_re_out(1214),
            data_re_in(63) => mul_re_out(1215),
            data_im_in(0) => mul_im_out(1152),
            data_im_in(1) => mul_im_out(1153),
            data_im_in(2) => mul_im_out(1154),
            data_im_in(3) => mul_im_out(1155),
            data_im_in(4) => mul_im_out(1156),
            data_im_in(5) => mul_im_out(1157),
            data_im_in(6) => mul_im_out(1158),
            data_im_in(7) => mul_im_out(1159),
            data_im_in(8) => mul_im_out(1160),
            data_im_in(9) => mul_im_out(1161),
            data_im_in(10) => mul_im_out(1162),
            data_im_in(11) => mul_im_out(1163),
            data_im_in(12) => mul_im_out(1164),
            data_im_in(13) => mul_im_out(1165),
            data_im_in(14) => mul_im_out(1166),
            data_im_in(15) => mul_im_out(1167),
            data_im_in(16) => mul_im_out(1168),
            data_im_in(17) => mul_im_out(1169),
            data_im_in(18) => mul_im_out(1170),
            data_im_in(19) => mul_im_out(1171),
            data_im_in(20) => mul_im_out(1172),
            data_im_in(21) => mul_im_out(1173),
            data_im_in(22) => mul_im_out(1174),
            data_im_in(23) => mul_im_out(1175),
            data_im_in(24) => mul_im_out(1176),
            data_im_in(25) => mul_im_out(1177),
            data_im_in(26) => mul_im_out(1178),
            data_im_in(27) => mul_im_out(1179),
            data_im_in(28) => mul_im_out(1180),
            data_im_in(29) => mul_im_out(1181),
            data_im_in(30) => mul_im_out(1182),
            data_im_in(31) => mul_im_out(1183),
            data_im_in(32) => mul_im_out(1184),
            data_im_in(33) => mul_im_out(1185),
            data_im_in(34) => mul_im_out(1186),
            data_im_in(35) => mul_im_out(1187),
            data_im_in(36) => mul_im_out(1188),
            data_im_in(37) => mul_im_out(1189),
            data_im_in(38) => mul_im_out(1190),
            data_im_in(39) => mul_im_out(1191),
            data_im_in(40) => mul_im_out(1192),
            data_im_in(41) => mul_im_out(1193),
            data_im_in(42) => mul_im_out(1194),
            data_im_in(43) => mul_im_out(1195),
            data_im_in(44) => mul_im_out(1196),
            data_im_in(45) => mul_im_out(1197),
            data_im_in(46) => mul_im_out(1198),
            data_im_in(47) => mul_im_out(1199),
            data_im_in(48) => mul_im_out(1200),
            data_im_in(49) => mul_im_out(1201),
            data_im_in(50) => mul_im_out(1202),
            data_im_in(51) => mul_im_out(1203),
            data_im_in(52) => mul_im_out(1204),
            data_im_in(53) => mul_im_out(1205),
            data_im_in(54) => mul_im_out(1206),
            data_im_in(55) => mul_im_out(1207),
            data_im_in(56) => mul_im_out(1208),
            data_im_in(57) => mul_im_out(1209),
            data_im_in(58) => mul_im_out(1210),
            data_im_in(59) => mul_im_out(1211),
            data_im_in(60) => mul_im_out(1212),
            data_im_in(61) => mul_im_out(1213),
            data_im_in(62) => mul_im_out(1214),
            data_im_in(63) => mul_im_out(1215),
            data_re_out(0) => data_re_out(18),
            data_re_out(1) => data_re_out(50),
            data_re_out(2) => data_re_out(82),
            data_re_out(3) => data_re_out(114),
            data_re_out(4) => data_re_out(146),
            data_re_out(5) => data_re_out(178),
            data_re_out(6) => data_re_out(210),
            data_re_out(7) => data_re_out(242),
            data_re_out(8) => data_re_out(274),
            data_re_out(9) => data_re_out(306),
            data_re_out(10) => data_re_out(338),
            data_re_out(11) => data_re_out(370),
            data_re_out(12) => data_re_out(402),
            data_re_out(13) => data_re_out(434),
            data_re_out(14) => data_re_out(466),
            data_re_out(15) => data_re_out(498),
            data_re_out(16) => data_re_out(530),
            data_re_out(17) => data_re_out(562),
            data_re_out(18) => data_re_out(594),
            data_re_out(19) => data_re_out(626),
            data_re_out(20) => data_re_out(658),
            data_re_out(21) => data_re_out(690),
            data_re_out(22) => data_re_out(722),
            data_re_out(23) => data_re_out(754),
            data_re_out(24) => data_re_out(786),
            data_re_out(25) => data_re_out(818),
            data_re_out(26) => data_re_out(850),
            data_re_out(27) => data_re_out(882),
            data_re_out(28) => data_re_out(914),
            data_re_out(29) => data_re_out(946),
            data_re_out(30) => data_re_out(978),
            data_re_out(31) => data_re_out(1010),
            data_re_out(32) => data_re_out(1042),
            data_re_out(33) => data_re_out(1074),
            data_re_out(34) => data_re_out(1106),
            data_re_out(35) => data_re_out(1138),
            data_re_out(36) => data_re_out(1170),
            data_re_out(37) => data_re_out(1202),
            data_re_out(38) => data_re_out(1234),
            data_re_out(39) => data_re_out(1266),
            data_re_out(40) => data_re_out(1298),
            data_re_out(41) => data_re_out(1330),
            data_re_out(42) => data_re_out(1362),
            data_re_out(43) => data_re_out(1394),
            data_re_out(44) => data_re_out(1426),
            data_re_out(45) => data_re_out(1458),
            data_re_out(46) => data_re_out(1490),
            data_re_out(47) => data_re_out(1522),
            data_re_out(48) => data_re_out(1554),
            data_re_out(49) => data_re_out(1586),
            data_re_out(50) => data_re_out(1618),
            data_re_out(51) => data_re_out(1650),
            data_re_out(52) => data_re_out(1682),
            data_re_out(53) => data_re_out(1714),
            data_re_out(54) => data_re_out(1746),
            data_re_out(55) => data_re_out(1778),
            data_re_out(56) => data_re_out(1810),
            data_re_out(57) => data_re_out(1842),
            data_re_out(58) => data_re_out(1874),
            data_re_out(59) => data_re_out(1906),
            data_re_out(60) => data_re_out(1938),
            data_re_out(61) => data_re_out(1970),
            data_re_out(62) => data_re_out(2002),
            data_re_out(63) => data_re_out(2034),
            data_im_out(0) => data_im_out(18),
            data_im_out(1) => data_im_out(50),
            data_im_out(2) => data_im_out(82),
            data_im_out(3) => data_im_out(114),
            data_im_out(4) => data_im_out(146),
            data_im_out(5) => data_im_out(178),
            data_im_out(6) => data_im_out(210),
            data_im_out(7) => data_im_out(242),
            data_im_out(8) => data_im_out(274),
            data_im_out(9) => data_im_out(306),
            data_im_out(10) => data_im_out(338),
            data_im_out(11) => data_im_out(370),
            data_im_out(12) => data_im_out(402),
            data_im_out(13) => data_im_out(434),
            data_im_out(14) => data_im_out(466),
            data_im_out(15) => data_im_out(498),
            data_im_out(16) => data_im_out(530),
            data_im_out(17) => data_im_out(562),
            data_im_out(18) => data_im_out(594),
            data_im_out(19) => data_im_out(626),
            data_im_out(20) => data_im_out(658),
            data_im_out(21) => data_im_out(690),
            data_im_out(22) => data_im_out(722),
            data_im_out(23) => data_im_out(754),
            data_im_out(24) => data_im_out(786),
            data_im_out(25) => data_im_out(818),
            data_im_out(26) => data_im_out(850),
            data_im_out(27) => data_im_out(882),
            data_im_out(28) => data_im_out(914),
            data_im_out(29) => data_im_out(946),
            data_im_out(30) => data_im_out(978),
            data_im_out(31) => data_im_out(1010),
            data_im_out(32) => data_im_out(1042),
            data_im_out(33) => data_im_out(1074),
            data_im_out(34) => data_im_out(1106),
            data_im_out(35) => data_im_out(1138),
            data_im_out(36) => data_im_out(1170),
            data_im_out(37) => data_im_out(1202),
            data_im_out(38) => data_im_out(1234),
            data_im_out(39) => data_im_out(1266),
            data_im_out(40) => data_im_out(1298),
            data_im_out(41) => data_im_out(1330),
            data_im_out(42) => data_im_out(1362),
            data_im_out(43) => data_im_out(1394),
            data_im_out(44) => data_im_out(1426),
            data_im_out(45) => data_im_out(1458),
            data_im_out(46) => data_im_out(1490),
            data_im_out(47) => data_im_out(1522),
            data_im_out(48) => data_im_out(1554),
            data_im_out(49) => data_im_out(1586),
            data_im_out(50) => data_im_out(1618),
            data_im_out(51) => data_im_out(1650),
            data_im_out(52) => data_im_out(1682),
            data_im_out(53) => data_im_out(1714),
            data_im_out(54) => data_im_out(1746),
            data_im_out(55) => data_im_out(1778),
            data_im_out(56) => data_im_out(1810),
            data_im_out(57) => data_im_out(1842),
            data_im_out(58) => data_im_out(1874),
            data_im_out(59) => data_im_out(1906),
            data_im_out(60) => data_im_out(1938),
            data_im_out(61) => data_im_out(1970),
            data_im_out(62) => data_im_out(2002),
            data_im_out(63) => data_im_out(2034)
        );           

    URFFT_PT64_19 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1216),
            data_re_in(1) => mul_re_out(1217),
            data_re_in(2) => mul_re_out(1218),
            data_re_in(3) => mul_re_out(1219),
            data_re_in(4) => mul_re_out(1220),
            data_re_in(5) => mul_re_out(1221),
            data_re_in(6) => mul_re_out(1222),
            data_re_in(7) => mul_re_out(1223),
            data_re_in(8) => mul_re_out(1224),
            data_re_in(9) => mul_re_out(1225),
            data_re_in(10) => mul_re_out(1226),
            data_re_in(11) => mul_re_out(1227),
            data_re_in(12) => mul_re_out(1228),
            data_re_in(13) => mul_re_out(1229),
            data_re_in(14) => mul_re_out(1230),
            data_re_in(15) => mul_re_out(1231),
            data_re_in(16) => mul_re_out(1232),
            data_re_in(17) => mul_re_out(1233),
            data_re_in(18) => mul_re_out(1234),
            data_re_in(19) => mul_re_out(1235),
            data_re_in(20) => mul_re_out(1236),
            data_re_in(21) => mul_re_out(1237),
            data_re_in(22) => mul_re_out(1238),
            data_re_in(23) => mul_re_out(1239),
            data_re_in(24) => mul_re_out(1240),
            data_re_in(25) => mul_re_out(1241),
            data_re_in(26) => mul_re_out(1242),
            data_re_in(27) => mul_re_out(1243),
            data_re_in(28) => mul_re_out(1244),
            data_re_in(29) => mul_re_out(1245),
            data_re_in(30) => mul_re_out(1246),
            data_re_in(31) => mul_re_out(1247),
            data_re_in(32) => mul_re_out(1248),
            data_re_in(33) => mul_re_out(1249),
            data_re_in(34) => mul_re_out(1250),
            data_re_in(35) => mul_re_out(1251),
            data_re_in(36) => mul_re_out(1252),
            data_re_in(37) => mul_re_out(1253),
            data_re_in(38) => mul_re_out(1254),
            data_re_in(39) => mul_re_out(1255),
            data_re_in(40) => mul_re_out(1256),
            data_re_in(41) => mul_re_out(1257),
            data_re_in(42) => mul_re_out(1258),
            data_re_in(43) => mul_re_out(1259),
            data_re_in(44) => mul_re_out(1260),
            data_re_in(45) => mul_re_out(1261),
            data_re_in(46) => mul_re_out(1262),
            data_re_in(47) => mul_re_out(1263),
            data_re_in(48) => mul_re_out(1264),
            data_re_in(49) => mul_re_out(1265),
            data_re_in(50) => mul_re_out(1266),
            data_re_in(51) => mul_re_out(1267),
            data_re_in(52) => mul_re_out(1268),
            data_re_in(53) => mul_re_out(1269),
            data_re_in(54) => mul_re_out(1270),
            data_re_in(55) => mul_re_out(1271),
            data_re_in(56) => mul_re_out(1272),
            data_re_in(57) => mul_re_out(1273),
            data_re_in(58) => mul_re_out(1274),
            data_re_in(59) => mul_re_out(1275),
            data_re_in(60) => mul_re_out(1276),
            data_re_in(61) => mul_re_out(1277),
            data_re_in(62) => mul_re_out(1278),
            data_re_in(63) => mul_re_out(1279),
            data_im_in(0) => mul_im_out(1216),
            data_im_in(1) => mul_im_out(1217),
            data_im_in(2) => mul_im_out(1218),
            data_im_in(3) => mul_im_out(1219),
            data_im_in(4) => mul_im_out(1220),
            data_im_in(5) => mul_im_out(1221),
            data_im_in(6) => mul_im_out(1222),
            data_im_in(7) => mul_im_out(1223),
            data_im_in(8) => mul_im_out(1224),
            data_im_in(9) => mul_im_out(1225),
            data_im_in(10) => mul_im_out(1226),
            data_im_in(11) => mul_im_out(1227),
            data_im_in(12) => mul_im_out(1228),
            data_im_in(13) => mul_im_out(1229),
            data_im_in(14) => mul_im_out(1230),
            data_im_in(15) => mul_im_out(1231),
            data_im_in(16) => mul_im_out(1232),
            data_im_in(17) => mul_im_out(1233),
            data_im_in(18) => mul_im_out(1234),
            data_im_in(19) => mul_im_out(1235),
            data_im_in(20) => mul_im_out(1236),
            data_im_in(21) => mul_im_out(1237),
            data_im_in(22) => mul_im_out(1238),
            data_im_in(23) => mul_im_out(1239),
            data_im_in(24) => mul_im_out(1240),
            data_im_in(25) => mul_im_out(1241),
            data_im_in(26) => mul_im_out(1242),
            data_im_in(27) => mul_im_out(1243),
            data_im_in(28) => mul_im_out(1244),
            data_im_in(29) => mul_im_out(1245),
            data_im_in(30) => mul_im_out(1246),
            data_im_in(31) => mul_im_out(1247),
            data_im_in(32) => mul_im_out(1248),
            data_im_in(33) => mul_im_out(1249),
            data_im_in(34) => mul_im_out(1250),
            data_im_in(35) => mul_im_out(1251),
            data_im_in(36) => mul_im_out(1252),
            data_im_in(37) => mul_im_out(1253),
            data_im_in(38) => mul_im_out(1254),
            data_im_in(39) => mul_im_out(1255),
            data_im_in(40) => mul_im_out(1256),
            data_im_in(41) => mul_im_out(1257),
            data_im_in(42) => mul_im_out(1258),
            data_im_in(43) => mul_im_out(1259),
            data_im_in(44) => mul_im_out(1260),
            data_im_in(45) => mul_im_out(1261),
            data_im_in(46) => mul_im_out(1262),
            data_im_in(47) => mul_im_out(1263),
            data_im_in(48) => mul_im_out(1264),
            data_im_in(49) => mul_im_out(1265),
            data_im_in(50) => mul_im_out(1266),
            data_im_in(51) => mul_im_out(1267),
            data_im_in(52) => mul_im_out(1268),
            data_im_in(53) => mul_im_out(1269),
            data_im_in(54) => mul_im_out(1270),
            data_im_in(55) => mul_im_out(1271),
            data_im_in(56) => mul_im_out(1272),
            data_im_in(57) => mul_im_out(1273),
            data_im_in(58) => mul_im_out(1274),
            data_im_in(59) => mul_im_out(1275),
            data_im_in(60) => mul_im_out(1276),
            data_im_in(61) => mul_im_out(1277),
            data_im_in(62) => mul_im_out(1278),
            data_im_in(63) => mul_im_out(1279),
            data_re_out(0) => data_re_out(19),
            data_re_out(1) => data_re_out(51),
            data_re_out(2) => data_re_out(83),
            data_re_out(3) => data_re_out(115),
            data_re_out(4) => data_re_out(147),
            data_re_out(5) => data_re_out(179),
            data_re_out(6) => data_re_out(211),
            data_re_out(7) => data_re_out(243),
            data_re_out(8) => data_re_out(275),
            data_re_out(9) => data_re_out(307),
            data_re_out(10) => data_re_out(339),
            data_re_out(11) => data_re_out(371),
            data_re_out(12) => data_re_out(403),
            data_re_out(13) => data_re_out(435),
            data_re_out(14) => data_re_out(467),
            data_re_out(15) => data_re_out(499),
            data_re_out(16) => data_re_out(531),
            data_re_out(17) => data_re_out(563),
            data_re_out(18) => data_re_out(595),
            data_re_out(19) => data_re_out(627),
            data_re_out(20) => data_re_out(659),
            data_re_out(21) => data_re_out(691),
            data_re_out(22) => data_re_out(723),
            data_re_out(23) => data_re_out(755),
            data_re_out(24) => data_re_out(787),
            data_re_out(25) => data_re_out(819),
            data_re_out(26) => data_re_out(851),
            data_re_out(27) => data_re_out(883),
            data_re_out(28) => data_re_out(915),
            data_re_out(29) => data_re_out(947),
            data_re_out(30) => data_re_out(979),
            data_re_out(31) => data_re_out(1011),
            data_re_out(32) => data_re_out(1043),
            data_re_out(33) => data_re_out(1075),
            data_re_out(34) => data_re_out(1107),
            data_re_out(35) => data_re_out(1139),
            data_re_out(36) => data_re_out(1171),
            data_re_out(37) => data_re_out(1203),
            data_re_out(38) => data_re_out(1235),
            data_re_out(39) => data_re_out(1267),
            data_re_out(40) => data_re_out(1299),
            data_re_out(41) => data_re_out(1331),
            data_re_out(42) => data_re_out(1363),
            data_re_out(43) => data_re_out(1395),
            data_re_out(44) => data_re_out(1427),
            data_re_out(45) => data_re_out(1459),
            data_re_out(46) => data_re_out(1491),
            data_re_out(47) => data_re_out(1523),
            data_re_out(48) => data_re_out(1555),
            data_re_out(49) => data_re_out(1587),
            data_re_out(50) => data_re_out(1619),
            data_re_out(51) => data_re_out(1651),
            data_re_out(52) => data_re_out(1683),
            data_re_out(53) => data_re_out(1715),
            data_re_out(54) => data_re_out(1747),
            data_re_out(55) => data_re_out(1779),
            data_re_out(56) => data_re_out(1811),
            data_re_out(57) => data_re_out(1843),
            data_re_out(58) => data_re_out(1875),
            data_re_out(59) => data_re_out(1907),
            data_re_out(60) => data_re_out(1939),
            data_re_out(61) => data_re_out(1971),
            data_re_out(62) => data_re_out(2003),
            data_re_out(63) => data_re_out(2035),
            data_im_out(0) => data_im_out(19),
            data_im_out(1) => data_im_out(51),
            data_im_out(2) => data_im_out(83),
            data_im_out(3) => data_im_out(115),
            data_im_out(4) => data_im_out(147),
            data_im_out(5) => data_im_out(179),
            data_im_out(6) => data_im_out(211),
            data_im_out(7) => data_im_out(243),
            data_im_out(8) => data_im_out(275),
            data_im_out(9) => data_im_out(307),
            data_im_out(10) => data_im_out(339),
            data_im_out(11) => data_im_out(371),
            data_im_out(12) => data_im_out(403),
            data_im_out(13) => data_im_out(435),
            data_im_out(14) => data_im_out(467),
            data_im_out(15) => data_im_out(499),
            data_im_out(16) => data_im_out(531),
            data_im_out(17) => data_im_out(563),
            data_im_out(18) => data_im_out(595),
            data_im_out(19) => data_im_out(627),
            data_im_out(20) => data_im_out(659),
            data_im_out(21) => data_im_out(691),
            data_im_out(22) => data_im_out(723),
            data_im_out(23) => data_im_out(755),
            data_im_out(24) => data_im_out(787),
            data_im_out(25) => data_im_out(819),
            data_im_out(26) => data_im_out(851),
            data_im_out(27) => data_im_out(883),
            data_im_out(28) => data_im_out(915),
            data_im_out(29) => data_im_out(947),
            data_im_out(30) => data_im_out(979),
            data_im_out(31) => data_im_out(1011),
            data_im_out(32) => data_im_out(1043),
            data_im_out(33) => data_im_out(1075),
            data_im_out(34) => data_im_out(1107),
            data_im_out(35) => data_im_out(1139),
            data_im_out(36) => data_im_out(1171),
            data_im_out(37) => data_im_out(1203),
            data_im_out(38) => data_im_out(1235),
            data_im_out(39) => data_im_out(1267),
            data_im_out(40) => data_im_out(1299),
            data_im_out(41) => data_im_out(1331),
            data_im_out(42) => data_im_out(1363),
            data_im_out(43) => data_im_out(1395),
            data_im_out(44) => data_im_out(1427),
            data_im_out(45) => data_im_out(1459),
            data_im_out(46) => data_im_out(1491),
            data_im_out(47) => data_im_out(1523),
            data_im_out(48) => data_im_out(1555),
            data_im_out(49) => data_im_out(1587),
            data_im_out(50) => data_im_out(1619),
            data_im_out(51) => data_im_out(1651),
            data_im_out(52) => data_im_out(1683),
            data_im_out(53) => data_im_out(1715),
            data_im_out(54) => data_im_out(1747),
            data_im_out(55) => data_im_out(1779),
            data_im_out(56) => data_im_out(1811),
            data_im_out(57) => data_im_out(1843),
            data_im_out(58) => data_im_out(1875),
            data_im_out(59) => data_im_out(1907),
            data_im_out(60) => data_im_out(1939),
            data_im_out(61) => data_im_out(1971),
            data_im_out(62) => data_im_out(2003),
            data_im_out(63) => data_im_out(2035)
        );           

    URFFT_PT64_20 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1280),
            data_re_in(1) => mul_re_out(1281),
            data_re_in(2) => mul_re_out(1282),
            data_re_in(3) => mul_re_out(1283),
            data_re_in(4) => mul_re_out(1284),
            data_re_in(5) => mul_re_out(1285),
            data_re_in(6) => mul_re_out(1286),
            data_re_in(7) => mul_re_out(1287),
            data_re_in(8) => mul_re_out(1288),
            data_re_in(9) => mul_re_out(1289),
            data_re_in(10) => mul_re_out(1290),
            data_re_in(11) => mul_re_out(1291),
            data_re_in(12) => mul_re_out(1292),
            data_re_in(13) => mul_re_out(1293),
            data_re_in(14) => mul_re_out(1294),
            data_re_in(15) => mul_re_out(1295),
            data_re_in(16) => mul_re_out(1296),
            data_re_in(17) => mul_re_out(1297),
            data_re_in(18) => mul_re_out(1298),
            data_re_in(19) => mul_re_out(1299),
            data_re_in(20) => mul_re_out(1300),
            data_re_in(21) => mul_re_out(1301),
            data_re_in(22) => mul_re_out(1302),
            data_re_in(23) => mul_re_out(1303),
            data_re_in(24) => mul_re_out(1304),
            data_re_in(25) => mul_re_out(1305),
            data_re_in(26) => mul_re_out(1306),
            data_re_in(27) => mul_re_out(1307),
            data_re_in(28) => mul_re_out(1308),
            data_re_in(29) => mul_re_out(1309),
            data_re_in(30) => mul_re_out(1310),
            data_re_in(31) => mul_re_out(1311),
            data_re_in(32) => mul_re_out(1312),
            data_re_in(33) => mul_re_out(1313),
            data_re_in(34) => mul_re_out(1314),
            data_re_in(35) => mul_re_out(1315),
            data_re_in(36) => mul_re_out(1316),
            data_re_in(37) => mul_re_out(1317),
            data_re_in(38) => mul_re_out(1318),
            data_re_in(39) => mul_re_out(1319),
            data_re_in(40) => mul_re_out(1320),
            data_re_in(41) => mul_re_out(1321),
            data_re_in(42) => mul_re_out(1322),
            data_re_in(43) => mul_re_out(1323),
            data_re_in(44) => mul_re_out(1324),
            data_re_in(45) => mul_re_out(1325),
            data_re_in(46) => mul_re_out(1326),
            data_re_in(47) => mul_re_out(1327),
            data_re_in(48) => mul_re_out(1328),
            data_re_in(49) => mul_re_out(1329),
            data_re_in(50) => mul_re_out(1330),
            data_re_in(51) => mul_re_out(1331),
            data_re_in(52) => mul_re_out(1332),
            data_re_in(53) => mul_re_out(1333),
            data_re_in(54) => mul_re_out(1334),
            data_re_in(55) => mul_re_out(1335),
            data_re_in(56) => mul_re_out(1336),
            data_re_in(57) => mul_re_out(1337),
            data_re_in(58) => mul_re_out(1338),
            data_re_in(59) => mul_re_out(1339),
            data_re_in(60) => mul_re_out(1340),
            data_re_in(61) => mul_re_out(1341),
            data_re_in(62) => mul_re_out(1342),
            data_re_in(63) => mul_re_out(1343),
            data_im_in(0) => mul_im_out(1280),
            data_im_in(1) => mul_im_out(1281),
            data_im_in(2) => mul_im_out(1282),
            data_im_in(3) => mul_im_out(1283),
            data_im_in(4) => mul_im_out(1284),
            data_im_in(5) => mul_im_out(1285),
            data_im_in(6) => mul_im_out(1286),
            data_im_in(7) => mul_im_out(1287),
            data_im_in(8) => mul_im_out(1288),
            data_im_in(9) => mul_im_out(1289),
            data_im_in(10) => mul_im_out(1290),
            data_im_in(11) => mul_im_out(1291),
            data_im_in(12) => mul_im_out(1292),
            data_im_in(13) => mul_im_out(1293),
            data_im_in(14) => mul_im_out(1294),
            data_im_in(15) => mul_im_out(1295),
            data_im_in(16) => mul_im_out(1296),
            data_im_in(17) => mul_im_out(1297),
            data_im_in(18) => mul_im_out(1298),
            data_im_in(19) => mul_im_out(1299),
            data_im_in(20) => mul_im_out(1300),
            data_im_in(21) => mul_im_out(1301),
            data_im_in(22) => mul_im_out(1302),
            data_im_in(23) => mul_im_out(1303),
            data_im_in(24) => mul_im_out(1304),
            data_im_in(25) => mul_im_out(1305),
            data_im_in(26) => mul_im_out(1306),
            data_im_in(27) => mul_im_out(1307),
            data_im_in(28) => mul_im_out(1308),
            data_im_in(29) => mul_im_out(1309),
            data_im_in(30) => mul_im_out(1310),
            data_im_in(31) => mul_im_out(1311),
            data_im_in(32) => mul_im_out(1312),
            data_im_in(33) => mul_im_out(1313),
            data_im_in(34) => mul_im_out(1314),
            data_im_in(35) => mul_im_out(1315),
            data_im_in(36) => mul_im_out(1316),
            data_im_in(37) => mul_im_out(1317),
            data_im_in(38) => mul_im_out(1318),
            data_im_in(39) => mul_im_out(1319),
            data_im_in(40) => mul_im_out(1320),
            data_im_in(41) => mul_im_out(1321),
            data_im_in(42) => mul_im_out(1322),
            data_im_in(43) => mul_im_out(1323),
            data_im_in(44) => mul_im_out(1324),
            data_im_in(45) => mul_im_out(1325),
            data_im_in(46) => mul_im_out(1326),
            data_im_in(47) => mul_im_out(1327),
            data_im_in(48) => mul_im_out(1328),
            data_im_in(49) => mul_im_out(1329),
            data_im_in(50) => mul_im_out(1330),
            data_im_in(51) => mul_im_out(1331),
            data_im_in(52) => mul_im_out(1332),
            data_im_in(53) => mul_im_out(1333),
            data_im_in(54) => mul_im_out(1334),
            data_im_in(55) => mul_im_out(1335),
            data_im_in(56) => mul_im_out(1336),
            data_im_in(57) => mul_im_out(1337),
            data_im_in(58) => mul_im_out(1338),
            data_im_in(59) => mul_im_out(1339),
            data_im_in(60) => mul_im_out(1340),
            data_im_in(61) => mul_im_out(1341),
            data_im_in(62) => mul_im_out(1342),
            data_im_in(63) => mul_im_out(1343),
            data_re_out(0) => data_re_out(20),
            data_re_out(1) => data_re_out(52),
            data_re_out(2) => data_re_out(84),
            data_re_out(3) => data_re_out(116),
            data_re_out(4) => data_re_out(148),
            data_re_out(5) => data_re_out(180),
            data_re_out(6) => data_re_out(212),
            data_re_out(7) => data_re_out(244),
            data_re_out(8) => data_re_out(276),
            data_re_out(9) => data_re_out(308),
            data_re_out(10) => data_re_out(340),
            data_re_out(11) => data_re_out(372),
            data_re_out(12) => data_re_out(404),
            data_re_out(13) => data_re_out(436),
            data_re_out(14) => data_re_out(468),
            data_re_out(15) => data_re_out(500),
            data_re_out(16) => data_re_out(532),
            data_re_out(17) => data_re_out(564),
            data_re_out(18) => data_re_out(596),
            data_re_out(19) => data_re_out(628),
            data_re_out(20) => data_re_out(660),
            data_re_out(21) => data_re_out(692),
            data_re_out(22) => data_re_out(724),
            data_re_out(23) => data_re_out(756),
            data_re_out(24) => data_re_out(788),
            data_re_out(25) => data_re_out(820),
            data_re_out(26) => data_re_out(852),
            data_re_out(27) => data_re_out(884),
            data_re_out(28) => data_re_out(916),
            data_re_out(29) => data_re_out(948),
            data_re_out(30) => data_re_out(980),
            data_re_out(31) => data_re_out(1012),
            data_re_out(32) => data_re_out(1044),
            data_re_out(33) => data_re_out(1076),
            data_re_out(34) => data_re_out(1108),
            data_re_out(35) => data_re_out(1140),
            data_re_out(36) => data_re_out(1172),
            data_re_out(37) => data_re_out(1204),
            data_re_out(38) => data_re_out(1236),
            data_re_out(39) => data_re_out(1268),
            data_re_out(40) => data_re_out(1300),
            data_re_out(41) => data_re_out(1332),
            data_re_out(42) => data_re_out(1364),
            data_re_out(43) => data_re_out(1396),
            data_re_out(44) => data_re_out(1428),
            data_re_out(45) => data_re_out(1460),
            data_re_out(46) => data_re_out(1492),
            data_re_out(47) => data_re_out(1524),
            data_re_out(48) => data_re_out(1556),
            data_re_out(49) => data_re_out(1588),
            data_re_out(50) => data_re_out(1620),
            data_re_out(51) => data_re_out(1652),
            data_re_out(52) => data_re_out(1684),
            data_re_out(53) => data_re_out(1716),
            data_re_out(54) => data_re_out(1748),
            data_re_out(55) => data_re_out(1780),
            data_re_out(56) => data_re_out(1812),
            data_re_out(57) => data_re_out(1844),
            data_re_out(58) => data_re_out(1876),
            data_re_out(59) => data_re_out(1908),
            data_re_out(60) => data_re_out(1940),
            data_re_out(61) => data_re_out(1972),
            data_re_out(62) => data_re_out(2004),
            data_re_out(63) => data_re_out(2036),
            data_im_out(0) => data_im_out(20),
            data_im_out(1) => data_im_out(52),
            data_im_out(2) => data_im_out(84),
            data_im_out(3) => data_im_out(116),
            data_im_out(4) => data_im_out(148),
            data_im_out(5) => data_im_out(180),
            data_im_out(6) => data_im_out(212),
            data_im_out(7) => data_im_out(244),
            data_im_out(8) => data_im_out(276),
            data_im_out(9) => data_im_out(308),
            data_im_out(10) => data_im_out(340),
            data_im_out(11) => data_im_out(372),
            data_im_out(12) => data_im_out(404),
            data_im_out(13) => data_im_out(436),
            data_im_out(14) => data_im_out(468),
            data_im_out(15) => data_im_out(500),
            data_im_out(16) => data_im_out(532),
            data_im_out(17) => data_im_out(564),
            data_im_out(18) => data_im_out(596),
            data_im_out(19) => data_im_out(628),
            data_im_out(20) => data_im_out(660),
            data_im_out(21) => data_im_out(692),
            data_im_out(22) => data_im_out(724),
            data_im_out(23) => data_im_out(756),
            data_im_out(24) => data_im_out(788),
            data_im_out(25) => data_im_out(820),
            data_im_out(26) => data_im_out(852),
            data_im_out(27) => data_im_out(884),
            data_im_out(28) => data_im_out(916),
            data_im_out(29) => data_im_out(948),
            data_im_out(30) => data_im_out(980),
            data_im_out(31) => data_im_out(1012),
            data_im_out(32) => data_im_out(1044),
            data_im_out(33) => data_im_out(1076),
            data_im_out(34) => data_im_out(1108),
            data_im_out(35) => data_im_out(1140),
            data_im_out(36) => data_im_out(1172),
            data_im_out(37) => data_im_out(1204),
            data_im_out(38) => data_im_out(1236),
            data_im_out(39) => data_im_out(1268),
            data_im_out(40) => data_im_out(1300),
            data_im_out(41) => data_im_out(1332),
            data_im_out(42) => data_im_out(1364),
            data_im_out(43) => data_im_out(1396),
            data_im_out(44) => data_im_out(1428),
            data_im_out(45) => data_im_out(1460),
            data_im_out(46) => data_im_out(1492),
            data_im_out(47) => data_im_out(1524),
            data_im_out(48) => data_im_out(1556),
            data_im_out(49) => data_im_out(1588),
            data_im_out(50) => data_im_out(1620),
            data_im_out(51) => data_im_out(1652),
            data_im_out(52) => data_im_out(1684),
            data_im_out(53) => data_im_out(1716),
            data_im_out(54) => data_im_out(1748),
            data_im_out(55) => data_im_out(1780),
            data_im_out(56) => data_im_out(1812),
            data_im_out(57) => data_im_out(1844),
            data_im_out(58) => data_im_out(1876),
            data_im_out(59) => data_im_out(1908),
            data_im_out(60) => data_im_out(1940),
            data_im_out(61) => data_im_out(1972),
            data_im_out(62) => data_im_out(2004),
            data_im_out(63) => data_im_out(2036)
        );           

    URFFT_PT64_21 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1344),
            data_re_in(1) => mul_re_out(1345),
            data_re_in(2) => mul_re_out(1346),
            data_re_in(3) => mul_re_out(1347),
            data_re_in(4) => mul_re_out(1348),
            data_re_in(5) => mul_re_out(1349),
            data_re_in(6) => mul_re_out(1350),
            data_re_in(7) => mul_re_out(1351),
            data_re_in(8) => mul_re_out(1352),
            data_re_in(9) => mul_re_out(1353),
            data_re_in(10) => mul_re_out(1354),
            data_re_in(11) => mul_re_out(1355),
            data_re_in(12) => mul_re_out(1356),
            data_re_in(13) => mul_re_out(1357),
            data_re_in(14) => mul_re_out(1358),
            data_re_in(15) => mul_re_out(1359),
            data_re_in(16) => mul_re_out(1360),
            data_re_in(17) => mul_re_out(1361),
            data_re_in(18) => mul_re_out(1362),
            data_re_in(19) => mul_re_out(1363),
            data_re_in(20) => mul_re_out(1364),
            data_re_in(21) => mul_re_out(1365),
            data_re_in(22) => mul_re_out(1366),
            data_re_in(23) => mul_re_out(1367),
            data_re_in(24) => mul_re_out(1368),
            data_re_in(25) => mul_re_out(1369),
            data_re_in(26) => mul_re_out(1370),
            data_re_in(27) => mul_re_out(1371),
            data_re_in(28) => mul_re_out(1372),
            data_re_in(29) => mul_re_out(1373),
            data_re_in(30) => mul_re_out(1374),
            data_re_in(31) => mul_re_out(1375),
            data_re_in(32) => mul_re_out(1376),
            data_re_in(33) => mul_re_out(1377),
            data_re_in(34) => mul_re_out(1378),
            data_re_in(35) => mul_re_out(1379),
            data_re_in(36) => mul_re_out(1380),
            data_re_in(37) => mul_re_out(1381),
            data_re_in(38) => mul_re_out(1382),
            data_re_in(39) => mul_re_out(1383),
            data_re_in(40) => mul_re_out(1384),
            data_re_in(41) => mul_re_out(1385),
            data_re_in(42) => mul_re_out(1386),
            data_re_in(43) => mul_re_out(1387),
            data_re_in(44) => mul_re_out(1388),
            data_re_in(45) => mul_re_out(1389),
            data_re_in(46) => mul_re_out(1390),
            data_re_in(47) => mul_re_out(1391),
            data_re_in(48) => mul_re_out(1392),
            data_re_in(49) => mul_re_out(1393),
            data_re_in(50) => mul_re_out(1394),
            data_re_in(51) => mul_re_out(1395),
            data_re_in(52) => mul_re_out(1396),
            data_re_in(53) => mul_re_out(1397),
            data_re_in(54) => mul_re_out(1398),
            data_re_in(55) => mul_re_out(1399),
            data_re_in(56) => mul_re_out(1400),
            data_re_in(57) => mul_re_out(1401),
            data_re_in(58) => mul_re_out(1402),
            data_re_in(59) => mul_re_out(1403),
            data_re_in(60) => mul_re_out(1404),
            data_re_in(61) => mul_re_out(1405),
            data_re_in(62) => mul_re_out(1406),
            data_re_in(63) => mul_re_out(1407),
            data_im_in(0) => mul_im_out(1344),
            data_im_in(1) => mul_im_out(1345),
            data_im_in(2) => mul_im_out(1346),
            data_im_in(3) => mul_im_out(1347),
            data_im_in(4) => mul_im_out(1348),
            data_im_in(5) => mul_im_out(1349),
            data_im_in(6) => mul_im_out(1350),
            data_im_in(7) => mul_im_out(1351),
            data_im_in(8) => mul_im_out(1352),
            data_im_in(9) => mul_im_out(1353),
            data_im_in(10) => mul_im_out(1354),
            data_im_in(11) => mul_im_out(1355),
            data_im_in(12) => mul_im_out(1356),
            data_im_in(13) => mul_im_out(1357),
            data_im_in(14) => mul_im_out(1358),
            data_im_in(15) => mul_im_out(1359),
            data_im_in(16) => mul_im_out(1360),
            data_im_in(17) => mul_im_out(1361),
            data_im_in(18) => mul_im_out(1362),
            data_im_in(19) => mul_im_out(1363),
            data_im_in(20) => mul_im_out(1364),
            data_im_in(21) => mul_im_out(1365),
            data_im_in(22) => mul_im_out(1366),
            data_im_in(23) => mul_im_out(1367),
            data_im_in(24) => mul_im_out(1368),
            data_im_in(25) => mul_im_out(1369),
            data_im_in(26) => mul_im_out(1370),
            data_im_in(27) => mul_im_out(1371),
            data_im_in(28) => mul_im_out(1372),
            data_im_in(29) => mul_im_out(1373),
            data_im_in(30) => mul_im_out(1374),
            data_im_in(31) => mul_im_out(1375),
            data_im_in(32) => mul_im_out(1376),
            data_im_in(33) => mul_im_out(1377),
            data_im_in(34) => mul_im_out(1378),
            data_im_in(35) => mul_im_out(1379),
            data_im_in(36) => mul_im_out(1380),
            data_im_in(37) => mul_im_out(1381),
            data_im_in(38) => mul_im_out(1382),
            data_im_in(39) => mul_im_out(1383),
            data_im_in(40) => mul_im_out(1384),
            data_im_in(41) => mul_im_out(1385),
            data_im_in(42) => mul_im_out(1386),
            data_im_in(43) => mul_im_out(1387),
            data_im_in(44) => mul_im_out(1388),
            data_im_in(45) => mul_im_out(1389),
            data_im_in(46) => mul_im_out(1390),
            data_im_in(47) => mul_im_out(1391),
            data_im_in(48) => mul_im_out(1392),
            data_im_in(49) => mul_im_out(1393),
            data_im_in(50) => mul_im_out(1394),
            data_im_in(51) => mul_im_out(1395),
            data_im_in(52) => mul_im_out(1396),
            data_im_in(53) => mul_im_out(1397),
            data_im_in(54) => mul_im_out(1398),
            data_im_in(55) => mul_im_out(1399),
            data_im_in(56) => mul_im_out(1400),
            data_im_in(57) => mul_im_out(1401),
            data_im_in(58) => mul_im_out(1402),
            data_im_in(59) => mul_im_out(1403),
            data_im_in(60) => mul_im_out(1404),
            data_im_in(61) => mul_im_out(1405),
            data_im_in(62) => mul_im_out(1406),
            data_im_in(63) => mul_im_out(1407),
            data_re_out(0) => data_re_out(21),
            data_re_out(1) => data_re_out(53),
            data_re_out(2) => data_re_out(85),
            data_re_out(3) => data_re_out(117),
            data_re_out(4) => data_re_out(149),
            data_re_out(5) => data_re_out(181),
            data_re_out(6) => data_re_out(213),
            data_re_out(7) => data_re_out(245),
            data_re_out(8) => data_re_out(277),
            data_re_out(9) => data_re_out(309),
            data_re_out(10) => data_re_out(341),
            data_re_out(11) => data_re_out(373),
            data_re_out(12) => data_re_out(405),
            data_re_out(13) => data_re_out(437),
            data_re_out(14) => data_re_out(469),
            data_re_out(15) => data_re_out(501),
            data_re_out(16) => data_re_out(533),
            data_re_out(17) => data_re_out(565),
            data_re_out(18) => data_re_out(597),
            data_re_out(19) => data_re_out(629),
            data_re_out(20) => data_re_out(661),
            data_re_out(21) => data_re_out(693),
            data_re_out(22) => data_re_out(725),
            data_re_out(23) => data_re_out(757),
            data_re_out(24) => data_re_out(789),
            data_re_out(25) => data_re_out(821),
            data_re_out(26) => data_re_out(853),
            data_re_out(27) => data_re_out(885),
            data_re_out(28) => data_re_out(917),
            data_re_out(29) => data_re_out(949),
            data_re_out(30) => data_re_out(981),
            data_re_out(31) => data_re_out(1013),
            data_re_out(32) => data_re_out(1045),
            data_re_out(33) => data_re_out(1077),
            data_re_out(34) => data_re_out(1109),
            data_re_out(35) => data_re_out(1141),
            data_re_out(36) => data_re_out(1173),
            data_re_out(37) => data_re_out(1205),
            data_re_out(38) => data_re_out(1237),
            data_re_out(39) => data_re_out(1269),
            data_re_out(40) => data_re_out(1301),
            data_re_out(41) => data_re_out(1333),
            data_re_out(42) => data_re_out(1365),
            data_re_out(43) => data_re_out(1397),
            data_re_out(44) => data_re_out(1429),
            data_re_out(45) => data_re_out(1461),
            data_re_out(46) => data_re_out(1493),
            data_re_out(47) => data_re_out(1525),
            data_re_out(48) => data_re_out(1557),
            data_re_out(49) => data_re_out(1589),
            data_re_out(50) => data_re_out(1621),
            data_re_out(51) => data_re_out(1653),
            data_re_out(52) => data_re_out(1685),
            data_re_out(53) => data_re_out(1717),
            data_re_out(54) => data_re_out(1749),
            data_re_out(55) => data_re_out(1781),
            data_re_out(56) => data_re_out(1813),
            data_re_out(57) => data_re_out(1845),
            data_re_out(58) => data_re_out(1877),
            data_re_out(59) => data_re_out(1909),
            data_re_out(60) => data_re_out(1941),
            data_re_out(61) => data_re_out(1973),
            data_re_out(62) => data_re_out(2005),
            data_re_out(63) => data_re_out(2037),
            data_im_out(0) => data_im_out(21),
            data_im_out(1) => data_im_out(53),
            data_im_out(2) => data_im_out(85),
            data_im_out(3) => data_im_out(117),
            data_im_out(4) => data_im_out(149),
            data_im_out(5) => data_im_out(181),
            data_im_out(6) => data_im_out(213),
            data_im_out(7) => data_im_out(245),
            data_im_out(8) => data_im_out(277),
            data_im_out(9) => data_im_out(309),
            data_im_out(10) => data_im_out(341),
            data_im_out(11) => data_im_out(373),
            data_im_out(12) => data_im_out(405),
            data_im_out(13) => data_im_out(437),
            data_im_out(14) => data_im_out(469),
            data_im_out(15) => data_im_out(501),
            data_im_out(16) => data_im_out(533),
            data_im_out(17) => data_im_out(565),
            data_im_out(18) => data_im_out(597),
            data_im_out(19) => data_im_out(629),
            data_im_out(20) => data_im_out(661),
            data_im_out(21) => data_im_out(693),
            data_im_out(22) => data_im_out(725),
            data_im_out(23) => data_im_out(757),
            data_im_out(24) => data_im_out(789),
            data_im_out(25) => data_im_out(821),
            data_im_out(26) => data_im_out(853),
            data_im_out(27) => data_im_out(885),
            data_im_out(28) => data_im_out(917),
            data_im_out(29) => data_im_out(949),
            data_im_out(30) => data_im_out(981),
            data_im_out(31) => data_im_out(1013),
            data_im_out(32) => data_im_out(1045),
            data_im_out(33) => data_im_out(1077),
            data_im_out(34) => data_im_out(1109),
            data_im_out(35) => data_im_out(1141),
            data_im_out(36) => data_im_out(1173),
            data_im_out(37) => data_im_out(1205),
            data_im_out(38) => data_im_out(1237),
            data_im_out(39) => data_im_out(1269),
            data_im_out(40) => data_im_out(1301),
            data_im_out(41) => data_im_out(1333),
            data_im_out(42) => data_im_out(1365),
            data_im_out(43) => data_im_out(1397),
            data_im_out(44) => data_im_out(1429),
            data_im_out(45) => data_im_out(1461),
            data_im_out(46) => data_im_out(1493),
            data_im_out(47) => data_im_out(1525),
            data_im_out(48) => data_im_out(1557),
            data_im_out(49) => data_im_out(1589),
            data_im_out(50) => data_im_out(1621),
            data_im_out(51) => data_im_out(1653),
            data_im_out(52) => data_im_out(1685),
            data_im_out(53) => data_im_out(1717),
            data_im_out(54) => data_im_out(1749),
            data_im_out(55) => data_im_out(1781),
            data_im_out(56) => data_im_out(1813),
            data_im_out(57) => data_im_out(1845),
            data_im_out(58) => data_im_out(1877),
            data_im_out(59) => data_im_out(1909),
            data_im_out(60) => data_im_out(1941),
            data_im_out(61) => data_im_out(1973),
            data_im_out(62) => data_im_out(2005),
            data_im_out(63) => data_im_out(2037)
        );           

    URFFT_PT64_22 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1408),
            data_re_in(1) => mul_re_out(1409),
            data_re_in(2) => mul_re_out(1410),
            data_re_in(3) => mul_re_out(1411),
            data_re_in(4) => mul_re_out(1412),
            data_re_in(5) => mul_re_out(1413),
            data_re_in(6) => mul_re_out(1414),
            data_re_in(7) => mul_re_out(1415),
            data_re_in(8) => mul_re_out(1416),
            data_re_in(9) => mul_re_out(1417),
            data_re_in(10) => mul_re_out(1418),
            data_re_in(11) => mul_re_out(1419),
            data_re_in(12) => mul_re_out(1420),
            data_re_in(13) => mul_re_out(1421),
            data_re_in(14) => mul_re_out(1422),
            data_re_in(15) => mul_re_out(1423),
            data_re_in(16) => mul_re_out(1424),
            data_re_in(17) => mul_re_out(1425),
            data_re_in(18) => mul_re_out(1426),
            data_re_in(19) => mul_re_out(1427),
            data_re_in(20) => mul_re_out(1428),
            data_re_in(21) => mul_re_out(1429),
            data_re_in(22) => mul_re_out(1430),
            data_re_in(23) => mul_re_out(1431),
            data_re_in(24) => mul_re_out(1432),
            data_re_in(25) => mul_re_out(1433),
            data_re_in(26) => mul_re_out(1434),
            data_re_in(27) => mul_re_out(1435),
            data_re_in(28) => mul_re_out(1436),
            data_re_in(29) => mul_re_out(1437),
            data_re_in(30) => mul_re_out(1438),
            data_re_in(31) => mul_re_out(1439),
            data_re_in(32) => mul_re_out(1440),
            data_re_in(33) => mul_re_out(1441),
            data_re_in(34) => mul_re_out(1442),
            data_re_in(35) => mul_re_out(1443),
            data_re_in(36) => mul_re_out(1444),
            data_re_in(37) => mul_re_out(1445),
            data_re_in(38) => mul_re_out(1446),
            data_re_in(39) => mul_re_out(1447),
            data_re_in(40) => mul_re_out(1448),
            data_re_in(41) => mul_re_out(1449),
            data_re_in(42) => mul_re_out(1450),
            data_re_in(43) => mul_re_out(1451),
            data_re_in(44) => mul_re_out(1452),
            data_re_in(45) => mul_re_out(1453),
            data_re_in(46) => mul_re_out(1454),
            data_re_in(47) => mul_re_out(1455),
            data_re_in(48) => mul_re_out(1456),
            data_re_in(49) => mul_re_out(1457),
            data_re_in(50) => mul_re_out(1458),
            data_re_in(51) => mul_re_out(1459),
            data_re_in(52) => mul_re_out(1460),
            data_re_in(53) => mul_re_out(1461),
            data_re_in(54) => mul_re_out(1462),
            data_re_in(55) => mul_re_out(1463),
            data_re_in(56) => mul_re_out(1464),
            data_re_in(57) => mul_re_out(1465),
            data_re_in(58) => mul_re_out(1466),
            data_re_in(59) => mul_re_out(1467),
            data_re_in(60) => mul_re_out(1468),
            data_re_in(61) => mul_re_out(1469),
            data_re_in(62) => mul_re_out(1470),
            data_re_in(63) => mul_re_out(1471),
            data_im_in(0) => mul_im_out(1408),
            data_im_in(1) => mul_im_out(1409),
            data_im_in(2) => mul_im_out(1410),
            data_im_in(3) => mul_im_out(1411),
            data_im_in(4) => mul_im_out(1412),
            data_im_in(5) => mul_im_out(1413),
            data_im_in(6) => mul_im_out(1414),
            data_im_in(7) => mul_im_out(1415),
            data_im_in(8) => mul_im_out(1416),
            data_im_in(9) => mul_im_out(1417),
            data_im_in(10) => mul_im_out(1418),
            data_im_in(11) => mul_im_out(1419),
            data_im_in(12) => mul_im_out(1420),
            data_im_in(13) => mul_im_out(1421),
            data_im_in(14) => mul_im_out(1422),
            data_im_in(15) => mul_im_out(1423),
            data_im_in(16) => mul_im_out(1424),
            data_im_in(17) => mul_im_out(1425),
            data_im_in(18) => mul_im_out(1426),
            data_im_in(19) => mul_im_out(1427),
            data_im_in(20) => mul_im_out(1428),
            data_im_in(21) => mul_im_out(1429),
            data_im_in(22) => mul_im_out(1430),
            data_im_in(23) => mul_im_out(1431),
            data_im_in(24) => mul_im_out(1432),
            data_im_in(25) => mul_im_out(1433),
            data_im_in(26) => mul_im_out(1434),
            data_im_in(27) => mul_im_out(1435),
            data_im_in(28) => mul_im_out(1436),
            data_im_in(29) => mul_im_out(1437),
            data_im_in(30) => mul_im_out(1438),
            data_im_in(31) => mul_im_out(1439),
            data_im_in(32) => mul_im_out(1440),
            data_im_in(33) => mul_im_out(1441),
            data_im_in(34) => mul_im_out(1442),
            data_im_in(35) => mul_im_out(1443),
            data_im_in(36) => mul_im_out(1444),
            data_im_in(37) => mul_im_out(1445),
            data_im_in(38) => mul_im_out(1446),
            data_im_in(39) => mul_im_out(1447),
            data_im_in(40) => mul_im_out(1448),
            data_im_in(41) => mul_im_out(1449),
            data_im_in(42) => mul_im_out(1450),
            data_im_in(43) => mul_im_out(1451),
            data_im_in(44) => mul_im_out(1452),
            data_im_in(45) => mul_im_out(1453),
            data_im_in(46) => mul_im_out(1454),
            data_im_in(47) => mul_im_out(1455),
            data_im_in(48) => mul_im_out(1456),
            data_im_in(49) => mul_im_out(1457),
            data_im_in(50) => mul_im_out(1458),
            data_im_in(51) => mul_im_out(1459),
            data_im_in(52) => mul_im_out(1460),
            data_im_in(53) => mul_im_out(1461),
            data_im_in(54) => mul_im_out(1462),
            data_im_in(55) => mul_im_out(1463),
            data_im_in(56) => mul_im_out(1464),
            data_im_in(57) => mul_im_out(1465),
            data_im_in(58) => mul_im_out(1466),
            data_im_in(59) => mul_im_out(1467),
            data_im_in(60) => mul_im_out(1468),
            data_im_in(61) => mul_im_out(1469),
            data_im_in(62) => mul_im_out(1470),
            data_im_in(63) => mul_im_out(1471),
            data_re_out(0) => data_re_out(22),
            data_re_out(1) => data_re_out(54),
            data_re_out(2) => data_re_out(86),
            data_re_out(3) => data_re_out(118),
            data_re_out(4) => data_re_out(150),
            data_re_out(5) => data_re_out(182),
            data_re_out(6) => data_re_out(214),
            data_re_out(7) => data_re_out(246),
            data_re_out(8) => data_re_out(278),
            data_re_out(9) => data_re_out(310),
            data_re_out(10) => data_re_out(342),
            data_re_out(11) => data_re_out(374),
            data_re_out(12) => data_re_out(406),
            data_re_out(13) => data_re_out(438),
            data_re_out(14) => data_re_out(470),
            data_re_out(15) => data_re_out(502),
            data_re_out(16) => data_re_out(534),
            data_re_out(17) => data_re_out(566),
            data_re_out(18) => data_re_out(598),
            data_re_out(19) => data_re_out(630),
            data_re_out(20) => data_re_out(662),
            data_re_out(21) => data_re_out(694),
            data_re_out(22) => data_re_out(726),
            data_re_out(23) => data_re_out(758),
            data_re_out(24) => data_re_out(790),
            data_re_out(25) => data_re_out(822),
            data_re_out(26) => data_re_out(854),
            data_re_out(27) => data_re_out(886),
            data_re_out(28) => data_re_out(918),
            data_re_out(29) => data_re_out(950),
            data_re_out(30) => data_re_out(982),
            data_re_out(31) => data_re_out(1014),
            data_re_out(32) => data_re_out(1046),
            data_re_out(33) => data_re_out(1078),
            data_re_out(34) => data_re_out(1110),
            data_re_out(35) => data_re_out(1142),
            data_re_out(36) => data_re_out(1174),
            data_re_out(37) => data_re_out(1206),
            data_re_out(38) => data_re_out(1238),
            data_re_out(39) => data_re_out(1270),
            data_re_out(40) => data_re_out(1302),
            data_re_out(41) => data_re_out(1334),
            data_re_out(42) => data_re_out(1366),
            data_re_out(43) => data_re_out(1398),
            data_re_out(44) => data_re_out(1430),
            data_re_out(45) => data_re_out(1462),
            data_re_out(46) => data_re_out(1494),
            data_re_out(47) => data_re_out(1526),
            data_re_out(48) => data_re_out(1558),
            data_re_out(49) => data_re_out(1590),
            data_re_out(50) => data_re_out(1622),
            data_re_out(51) => data_re_out(1654),
            data_re_out(52) => data_re_out(1686),
            data_re_out(53) => data_re_out(1718),
            data_re_out(54) => data_re_out(1750),
            data_re_out(55) => data_re_out(1782),
            data_re_out(56) => data_re_out(1814),
            data_re_out(57) => data_re_out(1846),
            data_re_out(58) => data_re_out(1878),
            data_re_out(59) => data_re_out(1910),
            data_re_out(60) => data_re_out(1942),
            data_re_out(61) => data_re_out(1974),
            data_re_out(62) => data_re_out(2006),
            data_re_out(63) => data_re_out(2038),
            data_im_out(0) => data_im_out(22),
            data_im_out(1) => data_im_out(54),
            data_im_out(2) => data_im_out(86),
            data_im_out(3) => data_im_out(118),
            data_im_out(4) => data_im_out(150),
            data_im_out(5) => data_im_out(182),
            data_im_out(6) => data_im_out(214),
            data_im_out(7) => data_im_out(246),
            data_im_out(8) => data_im_out(278),
            data_im_out(9) => data_im_out(310),
            data_im_out(10) => data_im_out(342),
            data_im_out(11) => data_im_out(374),
            data_im_out(12) => data_im_out(406),
            data_im_out(13) => data_im_out(438),
            data_im_out(14) => data_im_out(470),
            data_im_out(15) => data_im_out(502),
            data_im_out(16) => data_im_out(534),
            data_im_out(17) => data_im_out(566),
            data_im_out(18) => data_im_out(598),
            data_im_out(19) => data_im_out(630),
            data_im_out(20) => data_im_out(662),
            data_im_out(21) => data_im_out(694),
            data_im_out(22) => data_im_out(726),
            data_im_out(23) => data_im_out(758),
            data_im_out(24) => data_im_out(790),
            data_im_out(25) => data_im_out(822),
            data_im_out(26) => data_im_out(854),
            data_im_out(27) => data_im_out(886),
            data_im_out(28) => data_im_out(918),
            data_im_out(29) => data_im_out(950),
            data_im_out(30) => data_im_out(982),
            data_im_out(31) => data_im_out(1014),
            data_im_out(32) => data_im_out(1046),
            data_im_out(33) => data_im_out(1078),
            data_im_out(34) => data_im_out(1110),
            data_im_out(35) => data_im_out(1142),
            data_im_out(36) => data_im_out(1174),
            data_im_out(37) => data_im_out(1206),
            data_im_out(38) => data_im_out(1238),
            data_im_out(39) => data_im_out(1270),
            data_im_out(40) => data_im_out(1302),
            data_im_out(41) => data_im_out(1334),
            data_im_out(42) => data_im_out(1366),
            data_im_out(43) => data_im_out(1398),
            data_im_out(44) => data_im_out(1430),
            data_im_out(45) => data_im_out(1462),
            data_im_out(46) => data_im_out(1494),
            data_im_out(47) => data_im_out(1526),
            data_im_out(48) => data_im_out(1558),
            data_im_out(49) => data_im_out(1590),
            data_im_out(50) => data_im_out(1622),
            data_im_out(51) => data_im_out(1654),
            data_im_out(52) => data_im_out(1686),
            data_im_out(53) => data_im_out(1718),
            data_im_out(54) => data_im_out(1750),
            data_im_out(55) => data_im_out(1782),
            data_im_out(56) => data_im_out(1814),
            data_im_out(57) => data_im_out(1846),
            data_im_out(58) => data_im_out(1878),
            data_im_out(59) => data_im_out(1910),
            data_im_out(60) => data_im_out(1942),
            data_im_out(61) => data_im_out(1974),
            data_im_out(62) => data_im_out(2006),
            data_im_out(63) => data_im_out(2038)
        );           

    URFFT_PT64_23 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1472),
            data_re_in(1) => mul_re_out(1473),
            data_re_in(2) => mul_re_out(1474),
            data_re_in(3) => mul_re_out(1475),
            data_re_in(4) => mul_re_out(1476),
            data_re_in(5) => mul_re_out(1477),
            data_re_in(6) => mul_re_out(1478),
            data_re_in(7) => mul_re_out(1479),
            data_re_in(8) => mul_re_out(1480),
            data_re_in(9) => mul_re_out(1481),
            data_re_in(10) => mul_re_out(1482),
            data_re_in(11) => mul_re_out(1483),
            data_re_in(12) => mul_re_out(1484),
            data_re_in(13) => mul_re_out(1485),
            data_re_in(14) => mul_re_out(1486),
            data_re_in(15) => mul_re_out(1487),
            data_re_in(16) => mul_re_out(1488),
            data_re_in(17) => mul_re_out(1489),
            data_re_in(18) => mul_re_out(1490),
            data_re_in(19) => mul_re_out(1491),
            data_re_in(20) => mul_re_out(1492),
            data_re_in(21) => mul_re_out(1493),
            data_re_in(22) => mul_re_out(1494),
            data_re_in(23) => mul_re_out(1495),
            data_re_in(24) => mul_re_out(1496),
            data_re_in(25) => mul_re_out(1497),
            data_re_in(26) => mul_re_out(1498),
            data_re_in(27) => mul_re_out(1499),
            data_re_in(28) => mul_re_out(1500),
            data_re_in(29) => mul_re_out(1501),
            data_re_in(30) => mul_re_out(1502),
            data_re_in(31) => mul_re_out(1503),
            data_re_in(32) => mul_re_out(1504),
            data_re_in(33) => mul_re_out(1505),
            data_re_in(34) => mul_re_out(1506),
            data_re_in(35) => mul_re_out(1507),
            data_re_in(36) => mul_re_out(1508),
            data_re_in(37) => mul_re_out(1509),
            data_re_in(38) => mul_re_out(1510),
            data_re_in(39) => mul_re_out(1511),
            data_re_in(40) => mul_re_out(1512),
            data_re_in(41) => mul_re_out(1513),
            data_re_in(42) => mul_re_out(1514),
            data_re_in(43) => mul_re_out(1515),
            data_re_in(44) => mul_re_out(1516),
            data_re_in(45) => mul_re_out(1517),
            data_re_in(46) => mul_re_out(1518),
            data_re_in(47) => mul_re_out(1519),
            data_re_in(48) => mul_re_out(1520),
            data_re_in(49) => mul_re_out(1521),
            data_re_in(50) => mul_re_out(1522),
            data_re_in(51) => mul_re_out(1523),
            data_re_in(52) => mul_re_out(1524),
            data_re_in(53) => mul_re_out(1525),
            data_re_in(54) => mul_re_out(1526),
            data_re_in(55) => mul_re_out(1527),
            data_re_in(56) => mul_re_out(1528),
            data_re_in(57) => mul_re_out(1529),
            data_re_in(58) => mul_re_out(1530),
            data_re_in(59) => mul_re_out(1531),
            data_re_in(60) => mul_re_out(1532),
            data_re_in(61) => mul_re_out(1533),
            data_re_in(62) => mul_re_out(1534),
            data_re_in(63) => mul_re_out(1535),
            data_im_in(0) => mul_im_out(1472),
            data_im_in(1) => mul_im_out(1473),
            data_im_in(2) => mul_im_out(1474),
            data_im_in(3) => mul_im_out(1475),
            data_im_in(4) => mul_im_out(1476),
            data_im_in(5) => mul_im_out(1477),
            data_im_in(6) => mul_im_out(1478),
            data_im_in(7) => mul_im_out(1479),
            data_im_in(8) => mul_im_out(1480),
            data_im_in(9) => mul_im_out(1481),
            data_im_in(10) => mul_im_out(1482),
            data_im_in(11) => mul_im_out(1483),
            data_im_in(12) => mul_im_out(1484),
            data_im_in(13) => mul_im_out(1485),
            data_im_in(14) => mul_im_out(1486),
            data_im_in(15) => mul_im_out(1487),
            data_im_in(16) => mul_im_out(1488),
            data_im_in(17) => mul_im_out(1489),
            data_im_in(18) => mul_im_out(1490),
            data_im_in(19) => mul_im_out(1491),
            data_im_in(20) => mul_im_out(1492),
            data_im_in(21) => mul_im_out(1493),
            data_im_in(22) => mul_im_out(1494),
            data_im_in(23) => mul_im_out(1495),
            data_im_in(24) => mul_im_out(1496),
            data_im_in(25) => mul_im_out(1497),
            data_im_in(26) => mul_im_out(1498),
            data_im_in(27) => mul_im_out(1499),
            data_im_in(28) => mul_im_out(1500),
            data_im_in(29) => mul_im_out(1501),
            data_im_in(30) => mul_im_out(1502),
            data_im_in(31) => mul_im_out(1503),
            data_im_in(32) => mul_im_out(1504),
            data_im_in(33) => mul_im_out(1505),
            data_im_in(34) => mul_im_out(1506),
            data_im_in(35) => mul_im_out(1507),
            data_im_in(36) => mul_im_out(1508),
            data_im_in(37) => mul_im_out(1509),
            data_im_in(38) => mul_im_out(1510),
            data_im_in(39) => mul_im_out(1511),
            data_im_in(40) => mul_im_out(1512),
            data_im_in(41) => mul_im_out(1513),
            data_im_in(42) => mul_im_out(1514),
            data_im_in(43) => mul_im_out(1515),
            data_im_in(44) => mul_im_out(1516),
            data_im_in(45) => mul_im_out(1517),
            data_im_in(46) => mul_im_out(1518),
            data_im_in(47) => mul_im_out(1519),
            data_im_in(48) => mul_im_out(1520),
            data_im_in(49) => mul_im_out(1521),
            data_im_in(50) => mul_im_out(1522),
            data_im_in(51) => mul_im_out(1523),
            data_im_in(52) => mul_im_out(1524),
            data_im_in(53) => mul_im_out(1525),
            data_im_in(54) => mul_im_out(1526),
            data_im_in(55) => mul_im_out(1527),
            data_im_in(56) => mul_im_out(1528),
            data_im_in(57) => mul_im_out(1529),
            data_im_in(58) => mul_im_out(1530),
            data_im_in(59) => mul_im_out(1531),
            data_im_in(60) => mul_im_out(1532),
            data_im_in(61) => mul_im_out(1533),
            data_im_in(62) => mul_im_out(1534),
            data_im_in(63) => mul_im_out(1535),
            data_re_out(0) => data_re_out(23),
            data_re_out(1) => data_re_out(55),
            data_re_out(2) => data_re_out(87),
            data_re_out(3) => data_re_out(119),
            data_re_out(4) => data_re_out(151),
            data_re_out(5) => data_re_out(183),
            data_re_out(6) => data_re_out(215),
            data_re_out(7) => data_re_out(247),
            data_re_out(8) => data_re_out(279),
            data_re_out(9) => data_re_out(311),
            data_re_out(10) => data_re_out(343),
            data_re_out(11) => data_re_out(375),
            data_re_out(12) => data_re_out(407),
            data_re_out(13) => data_re_out(439),
            data_re_out(14) => data_re_out(471),
            data_re_out(15) => data_re_out(503),
            data_re_out(16) => data_re_out(535),
            data_re_out(17) => data_re_out(567),
            data_re_out(18) => data_re_out(599),
            data_re_out(19) => data_re_out(631),
            data_re_out(20) => data_re_out(663),
            data_re_out(21) => data_re_out(695),
            data_re_out(22) => data_re_out(727),
            data_re_out(23) => data_re_out(759),
            data_re_out(24) => data_re_out(791),
            data_re_out(25) => data_re_out(823),
            data_re_out(26) => data_re_out(855),
            data_re_out(27) => data_re_out(887),
            data_re_out(28) => data_re_out(919),
            data_re_out(29) => data_re_out(951),
            data_re_out(30) => data_re_out(983),
            data_re_out(31) => data_re_out(1015),
            data_re_out(32) => data_re_out(1047),
            data_re_out(33) => data_re_out(1079),
            data_re_out(34) => data_re_out(1111),
            data_re_out(35) => data_re_out(1143),
            data_re_out(36) => data_re_out(1175),
            data_re_out(37) => data_re_out(1207),
            data_re_out(38) => data_re_out(1239),
            data_re_out(39) => data_re_out(1271),
            data_re_out(40) => data_re_out(1303),
            data_re_out(41) => data_re_out(1335),
            data_re_out(42) => data_re_out(1367),
            data_re_out(43) => data_re_out(1399),
            data_re_out(44) => data_re_out(1431),
            data_re_out(45) => data_re_out(1463),
            data_re_out(46) => data_re_out(1495),
            data_re_out(47) => data_re_out(1527),
            data_re_out(48) => data_re_out(1559),
            data_re_out(49) => data_re_out(1591),
            data_re_out(50) => data_re_out(1623),
            data_re_out(51) => data_re_out(1655),
            data_re_out(52) => data_re_out(1687),
            data_re_out(53) => data_re_out(1719),
            data_re_out(54) => data_re_out(1751),
            data_re_out(55) => data_re_out(1783),
            data_re_out(56) => data_re_out(1815),
            data_re_out(57) => data_re_out(1847),
            data_re_out(58) => data_re_out(1879),
            data_re_out(59) => data_re_out(1911),
            data_re_out(60) => data_re_out(1943),
            data_re_out(61) => data_re_out(1975),
            data_re_out(62) => data_re_out(2007),
            data_re_out(63) => data_re_out(2039),
            data_im_out(0) => data_im_out(23),
            data_im_out(1) => data_im_out(55),
            data_im_out(2) => data_im_out(87),
            data_im_out(3) => data_im_out(119),
            data_im_out(4) => data_im_out(151),
            data_im_out(5) => data_im_out(183),
            data_im_out(6) => data_im_out(215),
            data_im_out(7) => data_im_out(247),
            data_im_out(8) => data_im_out(279),
            data_im_out(9) => data_im_out(311),
            data_im_out(10) => data_im_out(343),
            data_im_out(11) => data_im_out(375),
            data_im_out(12) => data_im_out(407),
            data_im_out(13) => data_im_out(439),
            data_im_out(14) => data_im_out(471),
            data_im_out(15) => data_im_out(503),
            data_im_out(16) => data_im_out(535),
            data_im_out(17) => data_im_out(567),
            data_im_out(18) => data_im_out(599),
            data_im_out(19) => data_im_out(631),
            data_im_out(20) => data_im_out(663),
            data_im_out(21) => data_im_out(695),
            data_im_out(22) => data_im_out(727),
            data_im_out(23) => data_im_out(759),
            data_im_out(24) => data_im_out(791),
            data_im_out(25) => data_im_out(823),
            data_im_out(26) => data_im_out(855),
            data_im_out(27) => data_im_out(887),
            data_im_out(28) => data_im_out(919),
            data_im_out(29) => data_im_out(951),
            data_im_out(30) => data_im_out(983),
            data_im_out(31) => data_im_out(1015),
            data_im_out(32) => data_im_out(1047),
            data_im_out(33) => data_im_out(1079),
            data_im_out(34) => data_im_out(1111),
            data_im_out(35) => data_im_out(1143),
            data_im_out(36) => data_im_out(1175),
            data_im_out(37) => data_im_out(1207),
            data_im_out(38) => data_im_out(1239),
            data_im_out(39) => data_im_out(1271),
            data_im_out(40) => data_im_out(1303),
            data_im_out(41) => data_im_out(1335),
            data_im_out(42) => data_im_out(1367),
            data_im_out(43) => data_im_out(1399),
            data_im_out(44) => data_im_out(1431),
            data_im_out(45) => data_im_out(1463),
            data_im_out(46) => data_im_out(1495),
            data_im_out(47) => data_im_out(1527),
            data_im_out(48) => data_im_out(1559),
            data_im_out(49) => data_im_out(1591),
            data_im_out(50) => data_im_out(1623),
            data_im_out(51) => data_im_out(1655),
            data_im_out(52) => data_im_out(1687),
            data_im_out(53) => data_im_out(1719),
            data_im_out(54) => data_im_out(1751),
            data_im_out(55) => data_im_out(1783),
            data_im_out(56) => data_im_out(1815),
            data_im_out(57) => data_im_out(1847),
            data_im_out(58) => data_im_out(1879),
            data_im_out(59) => data_im_out(1911),
            data_im_out(60) => data_im_out(1943),
            data_im_out(61) => data_im_out(1975),
            data_im_out(62) => data_im_out(2007),
            data_im_out(63) => data_im_out(2039)
        );           

    URFFT_PT64_24 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1536),
            data_re_in(1) => mul_re_out(1537),
            data_re_in(2) => mul_re_out(1538),
            data_re_in(3) => mul_re_out(1539),
            data_re_in(4) => mul_re_out(1540),
            data_re_in(5) => mul_re_out(1541),
            data_re_in(6) => mul_re_out(1542),
            data_re_in(7) => mul_re_out(1543),
            data_re_in(8) => mul_re_out(1544),
            data_re_in(9) => mul_re_out(1545),
            data_re_in(10) => mul_re_out(1546),
            data_re_in(11) => mul_re_out(1547),
            data_re_in(12) => mul_re_out(1548),
            data_re_in(13) => mul_re_out(1549),
            data_re_in(14) => mul_re_out(1550),
            data_re_in(15) => mul_re_out(1551),
            data_re_in(16) => mul_re_out(1552),
            data_re_in(17) => mul_re_out(1553),
            data_re_in(18) => mul_re_out(1554),
            data_re_in(19) => mul_re_out(1555),
            data_re_in(20) => mul_re_out(1556),
            data_re_in(21) => mul_re_out(1557),
            data_re_in(22) => mul_re_out(1558),
            data_re_in(23) => mul_re_out(1559),
            data_re_in(24) => mul_re_out(1560),
            data_re_in(25) => mul_re_out(1561),
            data_re_in(26) => mul_re_out(1562),
            data_re_in(27) => mul_re_out(1563),
            data_re_in(28) => mul_re_out(1564),
            data_re_in(29) => mul_re_out(1565),
            data_re_in(30) => mul_re_out(1566),
            data_re_in(31) => mul_re_out(1567),
            data_re_in(32) => mul_re_out(1568),
            data_re_in(33) => mul_re_out(1569),
            data_re_in(34) => mul_re_out(1570),
            data_re_in(35) => mul_re_out(1571),
            data_re_in(36) => mul_re_out(1572),
            data_re_in(37) => mul_re_out(1573),
            data_re_in(38) => mul_re_out(1574),
            data_re_in(39) => mul_re_out(1575),
            data_re_in(40) => mul_re_out(1576),
            data_re_in(41) => mul_re_out(1577),
            data_re_in(42) => mul_re_out(1578),
            data_re_in(43) => mul_re_out(1579),
            data_re_in(44) => mul_re_out(1580),
            data_re_in(45) => mul_re_out(1581),
            data_re_in(46) => mul_re_out(1582),
            data_re_in(47) => mul_re_out(1583),
            data_re_in(48) => mul_re_out(1584),
            data_re_in(49) => mul_re_out(1585),
            data_re_in(50) => mul_re_out(1586),
            data_re_in(51) => mul_re_out(1587),
            data_re_in(52) => mul_re_out(1588),
            data_re_in(53) => mul_re_out(1589),
            data_re_in(54) => mul_re_out(1590),
            data_re_in(55) => mul_re_out(1591),
            data_re_in(56) => mul_re_out(1592),
            data_re_in(57) => mul_re_out(1593),
            data_re_in(58) => mul_re_out(1594),
            data_re_in(59) => mul_re_out(1595),
            data_re_in(60) => mul_re_out(1596),
            data_re_in(61) => mul_re_out(1597),
            data_re_in(62) => mul_re_out(1598),
            data_re_in(63) => mul_re_out(1599),
            data_im_in(0) => mul_im_out(1536),
            data_im_in(1) => mul_im_out(1537),
            data_im_in(2) => mul_im_out(1538),
            data_im_in(3) => mul_im_out(1539),
            data_im_in(4) => mul_im_out(1540),
            data_im_in(5) => mul_im_out(1541),
            data_im_in(6) => mul_im_out(1542),
            data_im_in(7) => mul_im_out(1543),
            data_im_in(8) => mul_im_out(1544),
            data_im_in(9) => mul_im_out(1545),
            data_im_in(10) => mul_im_out(1546),
            data_im_in(11) => mul_im_out(1547),
            data_im_in(12) => mul_im_out(1548),
            data_im_in(13) => mul_im_out(1549),
            data_im_in(14) => mul_im_out(1550),
            data_im_in(15) => mul_im_out(1551),
            data_im_in(16) => mul_im_out(1552),
            data_im_in(17) => mul_im_out(1553),
            data_im_in(18) => mul_im_out(1554),
            data_im_in(19) => mul_im_out(1555),
            data_im_in(20) => mul_im_out(1556),
            data_im_in(21) => mul_im_out(1557),
            data_im_in(22) => mul_im_out(1558),
            data_im_in(23) => mul_im_out(1559),
            data_im_in(24) => mul_im_out(1560),
            data_im_in(25) => mul_im_out(1561),
            data_im_in(26) => mul_im_out(1562),
            data_im_in(27) => mul_im_out(1563),
            data_im_in(28) => mul_im_out(1564),
            data_im_in(29) => mul_im_out(1565),
            data_im_in(30) => mul_im_out(1566),
            data_im_in(31) => mul_im_out(1567),
            data_im_in(32) => mul_im_out(1568),
            data_im_in(33) => mul_im_out(1569),
            data_im_in(34) => mul_im_out(1570),
            data_im_in(35) => mul_im_out(1571),
            data_im_in(36) => mul_im_out(1572),
            data_im_in(37) => mul_im_out(1573),
            data_im_in(38) => mul_im_out(1574),
            data_im_in(39) => mul_im_out(1575),
            data_im_in(40) => mul_im_out(1576),
            data_im_in(41) => mul_im_out(1577),
            data_im_in(42) => mul_im_out(1578),
            data_im_in(43) => mul_im_out(1579),
            data_im_in(44) => mul_im_out(1580),
            data_im_in(45) => mul_im_out(1581),
            data_im_in(46) => mul_im_out(1582),
            data_im_in(47) => mul_im_out(1583),
            data_im_in(48) => mul_im_out(1584),
            data_im_in(49) => mul_im_out(1585),
            data_im_in(50) => mul_im_out(1586),
            data_im_in(51) => mul_im_out(1587),
            data_im_in(52) => mul_im_out(1588),
            data_im_in(53) => mul_im_out(1589),
            data_im_in(54) => mul_im_out(1590),
            data_im_in(55) => mul_im_out(1591),
            data_im_in(56) => mul_im_out(1592),
            data_im_in(57) => mul_im_out(1593),
            data_im_in(58) => mul_im_out(1594),
            data_im_in(59) => mul_im_out(1595),
            data_im_in(60) => mul_im_out(1596),
            data_im_in(61) => mul_im_out(1597),
            data_im_in(62) => mul_im_out(1598),
            data_im_in(63) => mul_im_out(1599),
            data_re_out(0) => data_re_out(24),
            data_re_out(1) => data_re_out(56),
            data_re_out(2) => data_re_out(88),
            data_re_out(3) => data_re_out(120),
            data_re_out(4) => data_re_out(152),
            data_re_out(5) => data_re_out(184),
            data_re_out(6) => data_re_out(216),
            data_re_out(7) => data_re_out(248),
            data_re_out(8) => data_re_out(280),
            data_re_out(9) => data_re_out(312),
            data_re_out(10) => data_re_out(344),
            data_re_out(11) => data_re_out(376),
            data_re_out(12) => data_re_out(408),
            data_re_out(13) => data_re_out(440),
            data_re_out(14) => data_re_out(472),
            data_re_out(15) => data_re_out(504),
            data_re_out(16) => data_re_out(536),
            data_re_out(17) => data_re_out(568),
            data_re_out(18) => data_re_out(600),
            data_re_out(19) => data_re_out(632),
            data_re_out(20) => data_re_out(664),
            data_re_out(21) => data_re_out(696),
            data_re_out(22) => data_re_out(728),
            data_re_out(23) => data_re_out(760),
            data_re_out(24) => data_re_out(792),
            data_re_out(25) => data_re_out(824),
            data_re_out(26) => data_re_out(856),
            data_re_out(27) => data_re_out(888),
            data_re_out(28) => data_re_out(920),
            data_re_out(29) => data_re_out(952),
            data_re_out(30) => data_re_out(984),
            data_re_out(31) => data_re_out(1016),
            data_re_out(32) => data_re_out(1048),
            data_re_out(33) => data_re_out(1080),
            data_re_out(34) => data_re_out(1112),
            data_re_out(35) => data_re_out(1144),
            data_re_out(36) => data_re_out(1176),
            data_re_out(37) => data_re_out(1208),
            data_re_out(38) => data_re_out(1240),
            data_re_out(39) => data_re_out(1272),
            data_re_out(40) => data_re_out(1304),
            data_re_out(41) => data_re_out(1336),
            data_re_out(42) => data_re_out(1368),
            data_re_out(43) => data_re_out(1400),
            data_re_out(44) => data_re_out(1432),
            data_re_out(45) => data_re_out(1464),
            data_re_out(46) => data_re_out(1496),
            data_re_out(47) => data_re_out(1528),
            data_re_out(48) => data_re_out(1560),
            data_re_out(49) => data_re_out(1592),
            data_re_out(50) => data_re_out(1624),
            data_re_out(51) => data_re_out(1656),
            data_re_out(52) => data_re_out(1688),
            data_re_out(53) => data_re_out(1720),
            data_re_out(54) => data_re_out(1752),
            data_re_out(55) => data_re_out(1784),
            data_re_out(56) => data_re_out(1816),
            data_re_out(57) => data_re_out(1848),
            data_re_out(58) => data_re_out(1880),
            data_re_out(59) => data_re_out(1912),
            data_re_out(60) => data_re_out(1944),
            data_re_out(61) => data_re_out(1976),
            data_re_out(62) => data_re_out(2008),
            data_re_out(63) => data_re_out(2040),
            data_im_out(0) => data_im_out(24),
            data_im_out(1) => data_im_out(56),
            data_im_out(2) => data_im_out(88),
            data_im_out(3) => data_im_out(120),
            data_im_out(4) => data_im_out(152),
            data_im_out(5) => data_im_out(184),
            data_im_out(6) => data_im_out(216),
            data_im_out(7) => data_im_out(248),
            data_im_out(8) => data_im_out(280),
            data_im_out(9) => data_im_out(312),
            data_im_out(10) => data_im_out(344),
            data_im_out(11) => data_im_out(376),
            data_im_out(12) => data_im_out(408),
            data_im_out(13) => data_im_out(440),
            data_im_out(14) => data_im_out(472),
            data_im_out(15) => data_im_out(504),
            data_im_out(16) => data_im_out(536),
            data_im_out(17) => data_im_out(568),
            data_im_out(18) => data_im_out(600),
            data_im_out(19) => data_im_out(632),
            data_im_out(20) => data_im_out(664),
            data_im_out(21) => data_im_out(696),
            data_im_out(22) => data_im_out(728),
            data_im_out(23) => data_im_out(760),
            data_im_out(24) => data_im_out(792),
            data_im_out(25) => data_im_out(824),
            data_im_out(26) => data_im_out(856),
            data_im_out(27) => data_im_out(888),
            data_im_out(28) => data_im_out(920),
            data_im_out(29) => data_im_out(952),
            data_im_out(30) => data_im_out(984),
            data_im_out(31) => data_im_out(1016),
            data_im_out(32) => data_im_out(1048),
            data_im_out(33) => data_im_out(1080),
            data_im_out(34) => data_im_out(1112),
            data_im_out(35) => data_im_out(1144),
            data_im_out(36) => data_im_out(1176),
            data_im_out(37) => data_im_out(1208),
            data_im_out(38) => data_im_out(1240),
            data_im_out(39) => data_im_out(1272),
            data_im_out(40) => data_im_out(1304),
            data_im_out(41) => data_im_out(1336),
            data_im_out(42) => data_im_out(1368),
            data_im_out(43) => data_im_out(1400),
            data_im_out(44) => data_im_out(1432),
            data_im_out(45) => data_im_out(1464),
            data_im_out(46) => data_im_out(1496),
            data_im_out(47) => data_im_out(1528),
            data_im_out(48) => data_im_out(1560),
            data_im_out(49) => data_im_out(1592),
            data_im_out(50) => data_im_out(1624),
            data_im_out(51) => data_im_out(1656),
            data_im_out(52) => data_im_out(1688),
            data_im_out(53) => data_im_out(1720),
            data_im_out(54) => data_im_out(1752),
            data_im_out(55) => data_im_out(1784),
            data_im_out(56) => data_im_out(1816),
            data_im_out(57) => data_im_out(1848),
            data_im_out(58) => data_im_out(1880),
            data_im_out(59) => data_im_out(1912),
            data_im_out(60) => data_im_out(1944),
            data_im_out(61) => data_im_out(1976),
            data_im_out(62) => data_im_out(2008),
            data_im_out(63) => data_im_out(2040)
        );           

    URFFT_PT64_25 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1600),
            data_re_in(1) => mul_re_out(1601),
            data_re_in(2) => mul_re_out(1602),
            data_re_in(3) => mul_re_out(1603),
            data_re_in(4) => mul_re_out(1604),
            data_re_in(5) => mul_re_out(1605),
            data_re_in(6) => mul_re_out(1606),
            data_re_in(7) => mul_re_out(1607),
            data_re_in(8) => mul_re_out(1608),
            data_re_in(9) => mul_re_out(1609),
            data_re_in(10) => mul_re_out(1610),
            data_re_in(11) => mul_re_out(1611),
            data_re_in(12) => mul_re_out(1612),
            data_re_in(13) => mul_re_out(1613),
            data_re_in(14) => mul_re_out(1614),
            data_re_in(15) => mul_re_out(1615),
            data_re_in(16) => mul_re_out(1616),
            data_re_in(17) => mul_re_out(1617),
            data_re_in(18) => mul_re_out(1618),
            data_re_in(19) => mul_re_out(1619),
            data_re_in(20) => mul_re_out(1620),
            data_re_in(21) => mul_re_out(1621),
            data_re_in(22) => mul_re_out(1622),
            data_re_in(23) => mul_re_out(1623),
            data_re_in(24) => mul_re_out(1624),
            data_re_in(25) => mul_re_out(1625),
            data_re_in(26) => mul_re_out(1626),
            data_re_in(27) => mul_re_out(1627),
            data_re_in(28) => mul_re_out(1628),
            data_re_in(29) => mul_re_out(1629),
            data_re_in(30) => mul_re_out(1630),
            data_re_in(31) => mul_re_out(1631),
            data_re_in(32) => mul_re_out(1632),
            data_re_in(33) => mul_re_out(1633),
            data_re_in(34) => mul_re_out(1634),
            data_re_in(35) => mul_re_out(1635),
            data_re_in(36) => mul_re_out(1636),
            data_re_in(37) => mul_re_out(1637),
            data_re_in(38) => mul_re_out(1638),
            data_re_in(39) => mul_re_out(1639),
            data_re_in(40) => mul_re_out(1640),
            data_re_in(41) => mul_re_out(1641),
            data_re_in(42) => mul_re_out(1642),
            data_re_in(43) => mul_re_out(1643),
            data_re_in(44) => mul_re_out(1644),
            data_re_in(45) => mul_re_out(1645),
            data_re_in(46) => mul_re_out(1646),
            data_re_in(47) => mul_re_out(1647),
            data_re_in(48) => mul_re_out(1648),
            data_re_in(49) => mul_re_out(1649),
            data_re_in(50) => mul_re_out(1650),
            data_re_in(51) => mul_re_out(1651),
            data_re_in(52) => mul_re_out(1652),
            data_re_in(53) => mul_re_out(1653),
            data_re_in(54) => mul_re_out(1654),
            data_re_in(55) => mul_re_out(1655),
            data_re_in(56) => mul_re_out(1656),
            data_re_in(57) => mul_re_out(1657),
            data_re_in(58) => mul_re_out(1658),
            data_re_in(59) => mul_re_out(1659),
            data_re_in(60) => mul_re_out(1660),
            data_re_in(61) => mul_re_out(1661),
            data_re_in(62) => mul_re_out(1662),
            data_re_in(63) => mul_re_out(1663),
            data_im_in(0) => mul_im_out(1600),
            data_im_in(1) => mul_im_out(1601),
            data_im_in(2) => mul_im_out(1602),
            data_im_in(3) => mul_im_out(1603),
            data_im_in(4) => mul_im_out(1604),
            data_im_in(5) => mul_im_out(1605),
            data_im_in(6) => mul_im_out(1606),
            data_im_in(7) => mul_im_out(1607),
            data_im_in(8) => mul_im_out(1608),
            data_im_in(9) => mul_im_out(1609),
            data_im_in(10) => mul_im_out(1610),
            data_im_in(11) => mul_im_out(1611),
            data_im_in(12) => mul_im_out(1612),
            data_im_in(13) => mul_im_out(1613),
            data_im_in(14) => mul_im_out(1614),
            data_im_in(15) => mul_im_out(1615),
            data_im_in(16) => mul_im_out(1616),
            data_im_in(17) => mul_im_out(1617),
            data_im_in(18) => mul_im_out(1618),
            data_im_in(19) => mul_im_out(1619),
            data_im_in(20) => mul_im_out(1620),
            data_im_in(21) => mul_im_out(1621),
            data_im_in(22) => mul_im_out(1622),
            data_im_in(23) => mul_im_out(1623),
            data_im_in(24) => mul_im_out(1624),
            data_im_in(25) => mul_im_out(1625),
            data_im_in(26) => mul_im_out(1626),
            data_im_in(27) => mul_im_out(1627),
            data_im_in(28) => mul_im_out(1628),
            data_im_in(29) => mul_im_out(1629),
            data_im_in(30) => mul_im_out(1630),
            data_im_in(31) => mul_im_out(1631),
            data_im_in(32) => mul_im_out(1632),
            data_im_in(33) => mul_im_out(1633),
            data_im_in(34) => mul_im_out(1634),
            data_im_in(35) => mul_im_out(1635),
            data_im_in(36) => mul_im_out(1636),
            data_im_in(37) => mul_im_out(1637),
            data_im_in(38) => mul_im_out(1638),
            data_im_in(39) => mul_im_out(1639),
            data_im_in(40) => mul_im_out(1640),
            data_im_in(41) => mul_im_out(1641),
            data_im_in(42) => mul_im_out(1642),
            data_im_in(43) => mul_im_out(1643),
            data_im_in(44) => mul_im_out(1644),
            data_im_in(45) => mul_im_out(1645),
            data_im_in(46) => mul_im_out(1646),
            data_im_in(47) => mul_im_out(1647),
            data_im_in(48) => mul_im_out(1648),
            data_im_in(49) => mul_im_out(1649),
            data_im_in(50) => mul_im_out(1650),
            data_im_in(51) => mul_im_out(1651),
            data_im_in(52) => mul_im_out(1652),
            data_im_in(53) => mul_im_out(1653),
            data_im_in(54) => mul_im_out(1654),
            data_im_in(55) => mul_im_out(1655),
            data_im_in(56) => mul_im_out(1656),
            data_im_in(57) => mul_im_out(1657),
            data_im_in(58) => mul_im_out(1658),
            data_im_in(59) => mul_im_out(1659),
            data_im_in(60) => mul_im_out(1660),
            data_im_in(61) => mul_im_out(1661),
            data_im_in(62) => mul_im_out(1662),
            data_im_in(63) => mul_im_out(1663),
            data_re_out(0) => data_re_out(25),
            data_re_out(1) => data_re_out(57),
            data_re_out(2) => data_re_out(89),
            data_re_out(3) => data_re_out(121),
            data_re_out(4) => data_re_out(153),
            data_re_out(5) => data_re_out(185),
            data_re_out(6) => data_re_out(217),
            data_re_out(7) => data_re_out(249),
            data_re_out(8) => data_re_out(281),
            data_re_out(9) => data_re_out(313),
            data_re_out(10) => data_re_out(345),
            data_re_out(11) => data_re_out(377),
            data_re_out(12) => data_re_out(409),
            data_re_out(13) => data_re_out(441),
            data_re_out(14) => data_re_out(473),
            data_re_out(15) => data_re_out(505),
            data_re_out(16) => data_re_out(537),
            data_re_out(17) => data_re_out(569),
            data_re_out(18) => data_re_out(601),
            data_re_out(19) => data_re_out(633),
            data_re_out(20) => data_re_out(665),
            data_re_out(21) => data_re_out(697),
            data_re_out(22) => data_re_out(729),
            data_re_out(23) => data_re_out(761),
            data_re_out(24) => data_re_out(793),
            data_re_out(25) => data_re_out(825),
            data_re_out(26) => data_re_out(857),
            data_re_out(27) => data_re_out(889),
            data_re_out(28) => data_re_out(921),
            data_re_out(29) => data_re_out(953),
            data_re_out(30) => data_re_out(985),
            data_re_out(31) => data_re_out(1017),
            data_re_out(32) => data_re_out(1049),
            data_re_out(33) => data_re_out(1081),
            data_re_out(34) => data_re_out(1113),
            data_re_out(35) => data_re_out(1145),
            data_re_out(36) => data_re_out(1177),
            data_re_out(37) => data_re_out(1209),
            data_re_out(38) => data_re_out(1241),
            data_re_out(39) => data_re_out(1273),
            data_re_out(40) => data_re_out(1305),
            data_re_out(41) => data_re_out(1337),
            data_re_out(42) => data_re_out(1369),
            data_re_out(43) => data_re_out(1401),
            data_re_out(44) => data_re_out(1433),
            data_re_out(45) => data_re_out(1465),
            data_re_out(46) => data_re_out(1497),
            data_re_out(47) => data_re_out(1529),
            data_re_out(48) => data_re_out(1561),
            data_re_out(49) => data_re_out(1593),
            data_re_out(50) => data_re_out(1625),
            data_re_out(51) => data_re_out(1657),
            data_re_out(52) => data_re_out(1689),
            data_re_out(53) => data_re_out(1721),
            data_re_out(54) => data_re_out(1753),
            data_re_out(55) => data_re_out(1785),
            data_re_out(56) => data_re_out(1817),
            data_re_out(57) => data_re_out(1849),
            data_re_out(58) => data_re_out(1881),
            data_re_out(59) => data_re_out(1913),
            data_re_out(60) => data_re_out(1945),
            data_re_out(61) => data_re_out(1977),
            data_re_out(62) => data_re_out(2009),
            data_re_out(63) => data_re_out(2041),
            data_im_out(0) => data_im_out(25),
            data_im_out(1) => data_im_out(57),
            data_im_out(2) => data_im_out(89),
            data_im_out(3) => data_im_out(121),
            data_im_out(4) => data_im_out(153),
            data_im_out(5) => data_im_out(185),
            data_im_out(6) => data_im_out(217),
            data_im_out(7) => data_im_out(249),
            data_im_out(8) => data_im_out(281),
            data_im_out(9) => data_im_out(313),
            data_im_out(10) => data_im_out(345),
            data_im_out(11) => data_im_out(377),
            data_im_out(12) => data_im_out(409),
            data_im_out(13) => data_im_out(441),
            data_im_out(14) => data_im_out(473),
            data_im_out(15) => data_im_out(505),
            data_im_out(16) => data_im_out(537),
            data_im_out(17) => data_im_out(569),
            data_im_out(18) => data_im_out(601),
            data_im_out(19) => data_im_out(633),
            data_im_out(20) => data_im_out(665),
            data_im_out(21) => data_im_out(697),
            data_im_out(22) => data_im_out(729),
            data_im_out(23) => data_im_out(761),
            data_im_out(24) => data_im_out(793),
            data_im_out(25) => data_im_out(825),
            data_im_out(26) => data_im_out(857),
            data_im_out(27) => data_im_out(889),
            data_im_out(28) => data_im_out(921),
            data_im_out(29) => data_im_out(953),
            data_im_out(30) => data_im_out(985),
            data_im_out(31) => data_im_out(1017),
            data_im_out(32) => data_im_out(1049),
            data_im_out(33) => data_im_out(1081),
            data_im_out(34) => data_im_out(1113),
            data_im_out(35) => data_im_out(1145),
            data_im_out(36) => data_im_out(1177),
            data_im_out(37) => data_im_out(1209),
            data_im_out(38) => data_im_out(1241),
            data_im_out(39) => data_im_out(1273),
            data_im_out(40) => data_im_out(1305),
            data_im_out(41) => data_im_out(1337),
            data_im_out(42) => data_im_out(1369),
            data_im_out(43) => data_im_out(1401),
            data_im_out(44) => data_im_out(1433),
            data_im_out(45) => data_im_out(1465),
            data_im_out(46) => data_im_out(1497),
            data_im_out(47) => data_im_out(1529),
            data_im_out(48) => data_im_out(1561),
            data_im_out(49) => data_im_out(1593),
            data_im_out(50) => data_im_out(1625),
            data_im_out(51) => data_im_out(1657),
            data_im_out(52) => data_im_out(1689),
            data_im_out(53) => data_im_out(1721),
            data_im_out(54) => data_im_out(1753),
            data_im_out(55) => data_im_out(1785),
            data_im_out(56) => data_im_out(1817),
            data_im_out(57) => data_im_out(1849),
            data_im_out(58) => data_im_out(1881),
            data_im_out(59) => data_im_out(1913),
            data_im_out(60) => data_im_out(1945),
            data_im_out(61) => data_im_out(1977),
            data_im_out(62) => data_im_out(2009),
            data_im_out(63) => data_im_out(2041)
        );           

    URFFT_PT64_26 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1664),
            data_re_in(1) => mul_re_out(1665),
            data_re_in(2) => mul_re_out(1666),
            data_re_in(3) => mul_re_out(1667),
            data_re_in(4) => mul_re_out(1668),
            data_re_in(5) => mul_re_out(1669),
            data_re_in(6) => mul_re_out(1670),
            data_re_in(7) => mul_re_out(1671),
            data_re_in(8) => mul_re_out(1672),
            data_re_in(9) => mul_re_out(1673),
            data_re_in(10) => mul_re_out(1674),
            data_re_in(11) => mul_re_out(1675),
            data_re_in(12) => mul_re_out(1676),
            data_re_in(13) => mul_re_out(1677),
            data_re_in(14) => mul_re_out(1678),
            data_re_in(15) => mul_re_out(1679),
            data_re_in(16) => mul_re_out(1680),
            data_re_in(17) => mul_re_out(1681),
            data_re_in(18) => mul_re_out(1682),
            data_re_in(19) => mul_re_out(1683),
            data_re_in(20) => mul_re_out(1684),
            data_re_in(21) => mul_re_out(1685),
            data_re_in(22) => mul_re_out(1686),
            data_re_in(23) => mul_re_out(1687),
            data_re_in(24) => mul_re_out(1688),
            data_re_in(25) => mul_re_out(1689),
            data_re_in(26) => mul_re_out(1690),
            data_re_in(27) => mul_re_out(1691),
            data_re_in(28) => mul_re_out(1692),
            data_re_in(29) => mul_re_out(1693),
            data_re_in(30) => mul_re_out(1694),
            data_re_in(31) => mul_re_out(1695),
            data_re_in(32) => mul_re_out(1696),
            data_re_in(33) => mul_re_out(1697),
            data_re_in(34) => mul_re_out(1698),
            data_re_in(35) => mul_re_out(1699),
            data_re_in(36) => mul_re_out(1700),
            data_re_in(37) => mul_re_out(1701),
            data_re_in(38) => mul_re_out(1702),
            data_re_in(39) => mul_re_out(1703),
            data_re_in(40) => mul_re_out(1704),
            data_re_in(41) => mul_re_out(1705),
            data_re_in(42) => mul_re_out(1706),
            data_re_in(43) => mul_re_out(1707),
            data_re_in(44) => mul_re_out(1708),
            data_re_in(45) => mul_re_out(1709),
            data_re_in(46) => mul_re_out(1710),
            data_re_in(47) => mul_re_out(1711),
            data_re_in(48) => mul_re_out(1712),
            data_re_in(49) => mul_re_out(1713),
            data_re_in(50) => mul_re_out(1714),
            data_re_in(51) => mul_re_out(1715),
            data_re_in(52) => mul_re_out(1716),
            data_re_in(53) => mul_re_out(1717),
            data_re_in(54) => mul_re_out(1718),
            data_re_in(55) => mul_re_out(1719),
            data_re_in(56) => mul_re_out(1720),
            data_re_in(57) => mul_re_out(1721),
            data_re_in(58) => mul_re_out(1722),
            data_re_in(59) => mul_re_out(1723),
            data_re_in(60) => mul_re_out(1724),
            data_re_in(61) => mul_re_out(1725),
            data_re_in(62) => mul_re_out(1726),
            data_re_in(63) => mul_re_out(1727),
            data_im_in(0) => mul_im_out(1664),
            data_im_in(1) => mul_im_out(1665),
            data_im_in(2) => mul_im_out(1666),
            data_im_in(3) => mul_im_out(1667),
            data_im_in(4) => mul_im_out(1668),
            data_im_in(5) => mul_im_out(1669),
            data_im_in(6) => mul_im_out(1670),
            data_im_in(7) => mul_im_out(1671),
            data_im_in(8) => mul_im_out(1672),
            data_im_in(9) => mul_im_out(1673),
            data_im_in(10) => mul_im_out(1674),
            data_im_in(11) => mul_im_out(1675),
            data_im_in(12) => mul_im_out(1676),
            data_im_in(13) => mul_im_out(1677),
            data_im_in(14) => mul_im_out(1678),
            data_im_in(15) => mul_im_out(1679),
            data_im_in(16) => mul_im_out(1680),
            data_im_in(17) => mul_im_out(1681),
            data_im_in(18) => mul_im_out(1682),
            data_im_in(19) => mul_im_out(1683),
            data_im_in(20) => mul_im_out(1684),
            data_im_in(21) => mul_im_out(1685),
            data_im_in(22) => mul_im_out(1686),
            data_im_in(23) => mul_im_out(1687),
            data_im_in(24) => mul_im_out(1688),
            data_im_in(25) => mul_im_out(1689),
            data_im_in(26) => mul_im_out(1690),
            data_im_in(27) => mul_im_out(1691),
            data_im_in(28) => mul_im_out(1692),
            data_im_in(29) => mul_im_out(1693),
            data_im_in(30) => mul_im_out(1694),
            data_im_in(31) => mul_im_out(1695),
            data_im_in(32) => mul_im_out(1696),
            data_im_in(33) => mul_im_out(1697),
            data_im_in(34) => mul_im_out(1698),
            data_im_in(35) => mul_im_out(1699),
            data_im_in(36) => mul_im_out(1700),
            data_im_in(37) => mul_im_out(1701),
            data_im_in(38) => mul_im_out(1702),
            data_im_in(39) => mul_im_out(1703),
            data_im_in(40) => mul_im_out(1704),
            data_im_in(41) => mul_im_out(1705),
            data_im_in(42) => mul_im_out(1706),
            data_im_in(43) => mul_im_out(1707),
            data_im_in(44) => mul_im_out(1708),
            data_im_in(45) => mul_im_out(1709),
            data_im_in(46) => mul_im_out(1710),
            data_im_in(47) => mul_im_out(1711),
            data_im_in(48) => mul_im_out(1712),
            data_im_in(49) => mul_im_out(1713),
            data_im_in(50) => mul_im_out(1714),
            data_im_in(51) => mul_im_out(1715),
            data_im_in(52) => mul_im_out(1716),
            data_im_in(53) => mul_im_out(1717),
            data_im_in(54) => mul_im_out(1718),
            data_im_in(55) => mul_im_out(1719),
            data_im_in(56) => mul_im_out(1720),
            data_im_in(57) => mul_im_out(1721),
            data_im_in(58) => mul_im_out(1722),
            data_im_in(59) => mul_im_out(1723),
            data_im_in(60) => mul_im_out(1724),
            data_im_in(61) => mul_im_out(1725),
            data_im_in(62) => mul_im_out(1726),
            data_im_in(63) => mul_im_out(1727),
            data_re_out(0) => data_re_out(26),
            data_re_out(1) => data_re_out(58),
            data_re_out(2) => data_re_out(90),
            data_re_out(3) => data_re_out(122),
            data_re_out(4) => data_re_out(154),
            data_re_out(5) => data_re_out(186),
            data_re_out(6) => data_re_out(218),
            data_re_out(7) => data_re_out(250),
            data_re_out(8) => data_re_out(282),
            data_re_out(9) => data_re_out(314),
            data_re_out(10) => data_re_out(346),
            data_re_out(11) => data_re_out(378),
            data_re_out(12) => data_re_out(410),
            data_re_out(13) => data_re_out(442),
            data_re_out(14) => data_re_out(474),
            data_re_out(15) => data_re_out(506),
            data_re_out(16) => data_re_out(538),
            data_re_out(17) => data_re_out(570),
            data_re_out(18) => data_re_out(602),
            data_re_out(19) => data_re_out(634),
            data_re_out(20) => data_re_out(666),
            data_re_out(21) => data_re_out(698),
            data_re_out(22) => data_re_out(730),
            data_re_out(23) => data_re_out(762),
            data_re_out(24) => data_re_out(794),
            data_re_out(25) => data_re_out(826),
            data_re_out(26) => data_re_out(858),
            data_re_out(27) => data_re_out(890),
            data_re_out(28) => data_re_out(922),
            data_re_out(29) => data_re_out(954),
            data_re_out(30) => data_re_out(986),
            data_re_out(31) => data_re_out(1018),
            data_re_out(32) => data_re_out(1050),
            data_re_out(33) => data_re_out(1082),
            data_re_out(34) => data_re_out(1114),
            data_re_out(35) => data_re_out(1146),
            data_re_out(36) => data_re_out(1178),
            data_re_out(37) => data_re_out(1210),
            data_re_out(38) => data_re_out(1242),
            data_re_out(39) => data_re_out(1274),
            data_re_out(40) => data_re_out(1306),
            data_re_out(41) => data_re_out(1338),
            data_re_out(42) => data_re_out(1370),
            data_re_out(43) => data_re_out(1402),
            data_re_out(44) => data_re_out(1434),
            data_re_out(45) => data_re_out(1466),
            data_re_out(46) => data_re_out(1498),
            data_re_out(47) => data_re_out(1530),
            data_re_out(48) => data_re_out(1562),
            data_re_out(49) => data_re_out(1594),
            data_re_out(50) => data_re_out(1626),
            data_re_out(51) => data_re_out(1658),
            data_re_out(52) => data_re_out(1690),
            data_re_out(53) => data_re_out(1722),
            data_re_out(54) => data_re_out(1754),
            data_re_out(55) => data_re_out(1786),
            data_re_out(56) => data_re_out(1818),
            data_re_out(57) => data_re_out(1850),
            data_re_out(58) => data_re_out(1882),
            data_re_out(59) => data_re_out(1914),
            data_re_out(60) => data_re_out(1946),
            data_re_out(61) => data_re_out(1978),
            data_re_out(62) => data_re_out(2010),
            data_re_out(63) => data_re_out(2042),
            data_im_out(0) => data_im_out(26),
            data_im_out(1) => data_im_out(58),
            data_im_out(2) => data_im_out(90),
            data_im_out(3) => data_im_out(122),
            data_im_out(4) => data_im_out(154),
            data_im_out(5) => data_im_out(186),
            data_im_out(6) => data_im_out(218),
            data_im_out(7) => data_im_out(250),
            data_im_out(8) => data_im_out(282),
            data_im_out(9) => data_im_out(314),
            data_im_out(10) => data_im_out(346),
            data_im_out(11) => data_im_out(378),
            data_im_out(12) => data_im_out(410),
            data_im_out(13) => data_im_out(442),
            data_im_out(14) => data_im_out(474),
            data_im_out(15) => data_im_out(506),
            data_im_out(16) => data_im_out(538),
            data_im_out(17) => data_im_out(570),
            data_im_out(18) => data_im_out(602),
            data_im_out(19) => data_im_out(634),
            data_im_out(20) => data_im_out(666),
            data_im_out(21) => data_im_out(698),
            data_im_out(22) => data_im_out(730),
            data_im_out(23) => data_im_out(762),
            data_im_out(24) => data_im_out(794),
            data_im_out(25) => data_im_out(826),
            data_im_out(26) => data_im_out(858),
            data_im_out(27) => data_im_out(890),
            data_im_out(28) => data_im_out(922),
            data_im_out(29) => data_im_out(954),
            data_im_out(30) => data_im_out(986),
            data_im_out(31) => data_im_out(1018),
            data_im_out(32) => data_im_out(1050),
            data_im_out(33) => data_im_out(1082),
            data_im_out(34) => data_im_out(1114),
            data_im_out(35) => data_im_out(1146),
            data_im_out(36) => data_im_out(1178),
            data_im_out(37) => data_im_out(1210),
            data_im_out(38) => data_im_out(1242),
            data_im_out(39) => data_im_out(1274),
            data_im_out(40) => data_im_out(1306),
            data_im_out(41) => data_im_out(1338),
            data_im_out(42) => data_im_out(1370),
            data_im_out(43) => data_im_out(1402),
            data_im_out(44) => data_im_out(1434),
            data_im_out(45) => data_im_out(1466),
            data_im_out(46) => data_im_out(1498),
            data_im_out(47) => data_im_out(1530),
            data_im_out(48) => data_im_out(1562),
            data_im_out(49) => data_im_out(1594),
            data_im_out(50) => data_im_out(1626),
            data_im_out(51) => data_im_out(1658),
            data_im_out(52) => data_im_out(1690),
            data_im_out(53) => data_im_out(1722),
            data_im_out(54) => data_im_out(1754),
            data_im_out(55) => data_im_out(1786),
            data_im_out(56) => data_im_out(1818),
            data_im_out(57) => data_im_out(1850),
            data_im_out(58) => data_im_out(1882),
            data_im_out(59) => data_im_out(1914),
            data_im_out(60) => data_im_out(1946),
            data_im_out(61) => data_im_out(1978),
            data_im_out(62) => data_im_out(2010),
            data_im_out(63) => data_im_out(2042)
        );           

    URFFT_PT64_27 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1728),
            data_re_in(1) => mul_re_out(1729),
            data_re_in(2) => mul_re_out(1730),
            data_re_in(3) => mul_re_out(1731),
            data_re_in(4) => mul_re_out(1732),
            data_re_in(5) => mul_re_out(1733),
            data_re_in(6) => mul_re_out(1734),
            data_re_in(7) => mul_re_out(1735),
            data_re_in(8) => mul_re_out(1736),
            data_re_in(9) => mul_re_out(1737),
            data_re_in(10) => mul_re_out(1738),
            data_re_in(11) => mul_re_out(1739),
            data_re_in(12) => mul_re_out(1740),
            data_re_in(13) => mul_re_out(1741),
            data_re_in(14) => mul_re_out(1742),
            data_re_in(15) => mul_re_out(1743),
            data_re_in(16) => mul_re_out(1744),
            data_re_in(17) => mul_re_out(1745),
            data_re_in(18) => mul_re_out(1746),
            data_re_in(19) => mul_re_out(1747),
            data_re_in(20) => mul_re_out(1748),
            data_re_in(21) => mul_re_out(1749),
            data_re_in(22) => mul_re_out(1750),
            data_re_in(23) => mul_re_out(1751),
            data_re_in(24) => mul_re_out(1752),
            data_re_in(25) => mul_re_out(1753),
            data_re_in(26) => mul_re_out(1754),
            data_re_in(27) => mul_re_out(1755),
            data_re_in(28) => mul_re_out(1756),
            data_re_in(29) => mul_re_out(1757),
            data_re_in(30) => mul_re_out(1758),
            data_re_in(31) => mul_re_out(1759),
            data_re_in(32) => mul_re_out(1760),
            data_re_in(33) => mul_re_out(1761),
            data_re_in(34) => mul_re_out(1762),
            data_re_in(35) => mul_re_out(1763),
            data_re_in(36) => mul_re_out(1764),
            data_re_in(37) => mul_re_out(1765),
            data_re_in(38) => mul_re_out(1766),
            data_re_in(39) => mul_re_out(1767),
            data_re_in(40) => mul_re_out(1768),
            data_re_in(41) => mul_re_out(1769),
            data_re_in(42) => mul_re_out(1770),
            data_re_in(43) => mul_re_out(1771),
            data_re_in(44) => mul_re_out(1772),
            data_re_in(45) => mul_re_out(1773),
            data_re_in(46) => mul_re_out(1774),
            data_re_in(47) => mul_re_out(1775),
            data_re_in(48) => mul_re_out(1776),
            data_re_in(49) => mul_re_out(1777),
            data_re_in(50) => mul_re_out(1778),
            data_re_in(51) => mul_re_out(1779),
            data_re_in(52) => mul_re_out(1780),
            data_re_in(53) => mul_re_out(1781),
            data_re_in(54) => mul_re_out(1782),
            data_re_in(55) => mul_re_out(1783),
            data_re_in(56) => mul_re_out(1784),
            data_re_in(57) => mul_re_out(1785),
            data_re_in(58) => mul_re_out(1786),
            data_re_in(59) => mul_re_out(1787),
            data_re_in(60) => mul_re_out(1788),
            data_re_in(61) => mul_re_out(1789),
            data_re_in(62) => mul_re_out(1790),
            data_re_in(63) => mul_re_out(1791),
            data_im_in(0) => mul_im_out(1728),
            data_im_in(1) => mul_im_out(1729),
            data_im_in(2) => mul_im_out(1730),
            data_im_in(3) => mul_im_out(1731),
            data_im_in(4) => mul_im_out(1732),
            data_im_in(5) => mul_im_out(1733),
            data_im_in(6) => mul_im_out(1734),
            data_im_in(7) => mul_im_out(1735),
            data_im_in(8) => mul_im_out(1736),
            data_im_in(9) => mul_im_out(1737),
            data_im_in(10) => mul_im_out(1738),
            data_im_in(11) => mul_im_out(1739),
            data_im_in(12) => mul_im_out(1740),
            data_im_in(13) => mul_im_out(1741),
            data_im_in(14) => mul_im_out(1742),
            data_im_in(15) => mul_im_out(1743),
            data_im_in(16) => mul_im_out(1744),
            data_im_in(17) => mul_im_out(1745),
            data_im_in(18) => mul_im_out(1746),
            data_im_in(19) => mul_im_out(1747),
            data_im_in(20) => mul_im_out(1748),
            data_im_in(21) => mul_im_out(1749),
            data_im_in(22) => mul_im_out(1750),
            data_im_in(23) => mul_im_out(1751),
            data_im_in(24) => mul_im_out(1752),
            data_im_in(25) => mul_im_out(1753),
            data_im_in(26) => mul_im_out(1754),
            data_im_in(27) => mul_im_out(1755),
            data_im_in(28) => mul_im_out(1756),
            data_im_in(29) => mul_im_out(1757),
            data_im_in(30) => mul_im_out(1758),
            data_im_in(31) => mul_im_out(1759),
            data_im_in(32) => mul_im_out(1760),
            data_im_in(33) => mul_im_out(1761),
            data_im_in(34) => mul_im_out(1762),
            data_im_in(35) => mul_im_out(1763),
            data_im_in(36) => mul_im_out(1764),
            data_im_in(37) => mul_im_out(1765),
            data_im_in(38) => mul_im_out(1766),
            data_im_in(39) => mul_im_out(1767),
            data_im_in(40) => mul_im_out(1768),
            data_im_in(41) => mul_im_out(1769),
            data_im_in(42) => mul_im_out(1770),
            data_im_in(43) => mul_im_out(1771),
            data_im_in(44) => mul_im_out(1772),
            data_im_in(45) => mul_im_out(1773),
            data_im_in(46) => mul_im_out(1774),
            data_im_in(47) => mul_im_out(1775),
            data_im_in(48) => mul_im_out(1776),
            data_im_in(49) => mul_im_out(1777),
            data_im_in(50) => mul_im_out(1778),
            data_im_in(51) => mul_im_out(1779),
            data_im_in(52) => mul_im_out(1780),
            data_im_in(53) => mul_im_out(1781),
            data_im_in(54) => mul_im_out(1782),
            data_im_in(55) => mul_im_out(1783),
            data_im_in(56) => mul_im_out(1784),
            data_im_in(57) => mul_im_out(1785),
            data_im_in(58) => mul_im_out(1786),
            data_im_in(59) => mul_im_out(1787),
            data_im_in(60) => mul_im_out(1788),
            data_im_in(61) => mul_im_out(1789),
            data_im_in(62) => mul_im_out(1790),
            data_im_in(63) => mul_im_out(1791),
            data_re_out(0) => data_re_out(27),
            data_re_out(1) => data_re_out(59),
            data_re_out(2) => data_re_out(91),
            data_re_out(3) => data_re_out(123),
            data_re_out(4) => data_re_out(155),
            data_re_out(5) => data_re_out(187),
            data_re_out(6) => data_re_out(219),
            data_re_out(7) => data_re_out(251),
            data_re_out(8) => data_re_out(283),
            data_re_out(9) => data_re_out(315),
            data_re_out(10) => data_re_out(347),
            data_re_out(11) => data_re_out(379),
            data_re_out(12) => data_re_out(411),
            data_re_out(13) => data_re_out(443),
            data_re_out(14) => data_re_out(475),
            data_re_out(15) => data_re_out(507),
            data_re_out(16) => data_re_out(539),
            data_re_out(17) => data_re_out(571),
            data_re_out(18) => data_re_out(603),
            data_re_out(19) => data_re_out(635),
            data_re_out(20) => data_re_out(667),
            data_re_out(21) => data_re_out(699),
            data_re_out(22) => data_re_out(731),
            data_re_out(23) => data_re_out(763),
            data_re_out(24) => data_re_out(795),
            data_re_out(25) => data_re_out(827),
            data_re_out(26) => data_re_out(859),
            data_re_out(27) => data_re_out(891),
            data_re_out(28) => data_re_out(923),
            data_re_out(29) => data_re_out(955),
            data_re_out(30) => data_re_out(987),
            data_re_out(31) => data_re_out(1019),
            data_re_out(32) => data_re_out(1051),
            data_re_out(33) => data_re_out(1083),
            data_re_out(34) => data_re_out(1115),
            data_re_out(35) => data_re_out(1147),
            data_re_out(36) => data_re_out(1179),
            data_re_out(37) => data_re_out(1211),
            data_re_out(38) => data_re_out(1243),
            data_re_out(39) => data_re_out(1275),
            data_re_out(40) => data_re_out(1307),
            data_re_out(41) => data_re_out(1339),
            data_re_out(42) => data_re_out(1371),
            data_re_out(43) => data_re_out(1403),
            data_re_out(44) => data_re_out(1435),
            data_re_out(45) => data_re_out(1467),
            data_re_out(46) => data_re_out(1499),
            data_re_out(47) => data_re_out(1531),
            data_re_out(48) => data_re_out(1563),
            data_re_out(49) => data_re_out(1595),
            data_re_out(50) => data_re_out(1627),
            data_re_out(51) => data_re_out(1659),
            data_re_out(52) => data_re_out(1691),
            data_re_out(53) => data_re_out(1723),
            data_re_out(54) => data_re_out(1755),
            data_re_out(55) => data_re_out(1787),
            data_re_out(56) => data_re_out(1819),
            data_re_out(57) => data_re_out(1851),
            data_re_out(58) => data_re_out(1883),
            data_re_out(59) => data_re_out(1915),
            data_re_out(60) => data_re_out(1947),
            data_re_out(61) => data_re_out(1979),
            data_re_out(62) => data_re_out(2011),
            data_re_out(63) => data_re_out(2043),
            data_im_out(0) => data_im_out(27),
            data_im_out(1) => data_im_out(59),
            data_im_out(2) => data_im_out(91),
            data_im_out(3) => data_im_out(123),
            data_im_out(4) => data_im_out(155),
            data_im_out(5) => data_im_out(187),
            data_im_out(6) => data_im_out(219),
            data_im_out(7) => data_im_out(251),
            data_im_out(8) => data_im_out(283),
            data_im_out(9) => data_im_out(315),
            data_im_out(10) => data_im_out(347),
            data_im_out(11) => data_im_out(379),
            data_im_out(12) => data_im_out(411),
            data_im_out(13) => data_im_out(443),
            data_im_out(14) => data_im_out(475),
            data_im_out(15) => data_im_out(507),
            data_im_out(16) => data_im_out(539),
            data_im_out(17) => data_im_out(571),
            data_im_out(18) => data_im_out(603),
            data_im_out(19) => data_im_out(635),
            data_im_out(20) => data_im_out(667),
            data_im_out(21) => data_im_out(699),
            data_im_out(22) => data_im_out(731),
            data_im_out(23) => data_im_out(763),
            data_im_out(24) => data_im_out(795),
            data_im_out(25) => data_im_out(827),
            data_im_out(26) => data_im_out(859),
            data_im_out(27) => data_im_out(891),
            data_im_out(28) => data_im_out(923),
            data_im_out(29) => data_im_out(955),
            data_im_out(30) => data_im_out(987),
            data_im_out(31) => data_im_out(1019),
            data_im_out(32) => data_im_out(1051),
            data_im_out(33) => data_im_out(1083),
            data_im_out(34) => data_im_out(1115),
            data_im_out(35) => data_im_out(1147),
            data_im_out(36) => data_im_out(1179),
            data_im_out(37) => data_im_out(1211),
            data_im_out(38) => data_im_out(1243),
            data_im_out(39) => data_im_out(1275),
            data_im_out(40) => data_im_out(1307),
            data_im_out(41) => data_im_out(1339),
            data_im_out(42) => data_im_out(1371),
            data_im_out(43) => data_im_out(1403),
            data_im_out(44) => data_im_out(1435),
            data_im_out(45) => data_im_out(1467),
            data_im_out(46) => data_im_out(1499),
            data_im_out(47) => data_im_out(1531),
            data_im_out(48) => data_im_out(1563),
            data_im_out(49) => data_im_out(1595),
            data_im_out(50) => data_im_out(1627),
            data_im_out(51) => data_im_out(1659),
            data_im_out(52) => data_im_out(1691),
            data_im_out(53) => data_im_out(1723),
            data_im_out(54) => data_im_out(1755),
            data_im_out(55) => data_im_out(1787),
            data_im_out(56) => data_im_out(1819),
            data_im_out(57) => data_im_out(1851),
            data_im_out(58) => data_im_out(1883),
            data_im_out(59) => data_im_out(1915),
            data_im_out(60) => data_im_out(1947),
            data_im_out(61) => data_im_out(1979),
            data_im_out(62) => data_im_out(2011),
            data_im_out(63) => data_im_out(2043)
        );           

    URFFT_PT64_28 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1792),
            data_re_in(1) => mul_re_out(1793),
            data_re_in(2) => mul_re_out(1794),
            data_re_in(3) => mul_re_out(1795),
            data_re_in(4) => mul_re_out(1796),
            data_re_in(5) => mul_re_out(1797),
            data_re_in(6) => mul_re_out(1798),
            data_re_in(7) => mul_re_out(1799),
            data_re_in(8) => mul_re_out(1800),
            data_re_in(9) => mul_re_out(1801),
            data_re_in(10) => mul_re_out(1802),
            data_re_in(11) => mul_re_out(1803),
            data_re_in(12) => mul_re_out(1804),
            data_re_in(13) => mul_re_out(1805),
            data_re_in(14) => mul_re_out(1806),
            data_re_in(15) => mul_re_out(1807),
            data_re_in(16) => mul_re_out(1808),
            data_re_in(17) => mul_re_out(1809),
            data_re_in(18) => mul_re_out(1810),
            data_re_in(19) => mul_re_out(1811),
            data_re_in(20) => mul_re_out(1812),
            data_re_in(21) => mul_re_out(1813),
            data_re_in(22) => mul_re_out(1814),
            data_re_in(23) => mul_re_out(1815),
            data_re_in(24) => mul_re_out(1816),
            data_re_in(25) => mul_re_out(1817),
            data_re_in(26) => mul_re_out(1818),
            data_re_in(27) => mul_re_out(1819),
            data_re_in(28) => mul_re_out(1820),
            data_re_in(29) => mul_re_out(1821),
            data_re_in(30) => mul_re_out(1822),
            data_re_in(31) => mul_re_out(1823),
            data_re_in(32) => mul_re_out(1824),
            data_re_in(33) => mul_re_out(1825),
            data_re_in(34) => mul_re_out(1826),
            data_re_in(35) => mul_re_out(1827),
            data_re_in(36) => mul_re_out(1828),
            data_re_in(37) => mul_re_out(1829),
            data_re_in(38) => mul_re_out(1830),
            data_re_in(39) => mul_re_out(1831),
            data_re_in(40) => mul_re_out(1832),
            data_re_in(41) => mul_re_out(1833),
            data_re_in(42) => mul_re_out(1834),
            data_re_in(43) => mul_re_out(1835),
            data_re_in(44) => mul_re_out(1836),
            data_re_in(45) => mul_re_out(1837),
            data_re_in(46) => mul_re_out(1838),
            data_re_in(47) => mul_re_out(1839),
            data_re_in(48) => mul_re_out(1840),
            data_re_in(49) => mul_re_out(1841),
            data_re_in(50) => mul_re_out(1842),
            data_re_in(51) => mul_re_out(1843),
            data_re_in(52) => mul_re_out(1844),
            data_re_in(53) => mul_re_out(1845),
            data_re_in(54) => mul_re_out(1846),
            data_re_in(55) => mul_re_out(1847),
            data_re_in(56) => mul_re_out(1848),
            data_re_in(57) => mul_re_out(1849),
            data_re_in(58) => mul_re_out(1850),
            data_re_in(59) => mul_re_out(1851),
            data_re_in(60) => mul_re_out(1852),
            data_re_in(61) => mul_re_out(1853),
            data_re_in(62) => mul_re_out(1854),
            data_re_in(63) => mul_re_out(1855),
            data_im_in(0) => mul_im_out(1792),
            data_im_in(1) => mul_im_out(1793),
            data_im_in(2) => mul_im_out(1794),
            data_im_in(3) => mul_im_out(1795),
            data_im_in(4) => mul_im_out(1796),
            data_im_in(5) => mul_im_out(1797),
            data_im_in(6) => mul_im_out(1798),
            data_im_in(7) => mul_im_out(1799),
            data_im_in(8) => mul_im_out(1800),
            data_im_in(9) => mul_im_out(1801),
            data_im_in(10) => mul_im_out(1802),
            data_im_in(11) => mul_im_out(1803),
            data_im_in(12) => mul_im_out(1804),
            data_im_in(13) => mul_im_out(1805),
            data_im_in(14) => mul_im_out(1806),
            data_im_in(15) => mul_im_out(1807),
            data_im_in(16) => mul_im_out(1808),
            data_im_in(17) => mul_im_out(1809),
            data_im_in(18) => mul_im_out(1810),
            data_im_in(19) => mul_im_out(1811),
            data_im_in(20) => mul_im_out(1812),
            data_im_in(21) => mul_im_out(1813),
            data_im_in(22) => mul_im_out(1814),
            data_im_in(23) => mul_im_out(1815),
            data_im_in(24) => mul_im_out(1816),
            data_im_in(25) => mul_im_out(1817),
            data_im_in(26) => mul_im_out(1818),
            data_im_in(27) => mul_im_out(1819),
            data_im_in(28) => mul_im_out(1820),
            data_im_in(29) => mul_im_out(1821),
            data_im_in(30) => mul_im_out(1822),
            data_im_in(31) => mul_im_out(1823),
            data_im_in(32) => mul_im_out(1824),
            data_im_in(33) => mul_im_out(1825),
            data_im_in(34) => mul_im_out(1826),
            data_im_in(35) => mul_im_out(1827),
            data_im_in(36) => mul_im_out(1828),
            data_im_in(37) => mul_im_out(1829),
            data_im_in(38) => mul_im_out(1830),
            data_im_in(39) => mul_im_out(1831),
            data_im_in(40) => mul_im_out(1832),
            data_im_in(41) => mul_im_out(1833),
            data_im_in(42) => mul_im_out(1834),
            data_im_in(43) => mul_im_out(1835),
            data_im_in(44) => mul_im_out(1836),
            data_im_in(45) => mul_im_out(1837),
            data_im_in(46) => mul_im_out(1838),
            data_im_in(47) => mul_im_out(1839),
            data_im_in(48) => mul_im_out(1840),
            data_im_in(49) => mul_im_out(1841),
            data_im_in(50) => mul_im_out(1842),
            data_im_in(51) => mul_im_out(1843),
            data_im_in(52) => mul_im_out(1844),
            data_im_in(53) => mul_im_out(1845),
            data_im_in(54) => mul_im_out(1846),
            data_im_in(55) => mul_im_out(1847),
            data_im_in(56) => mul_im_out(1848),
            data_im_in(57) => mul_im_out(1849),
            data_im_in(58) => mul_im_out(1850),
            data_im_in(59) => mul_im_out(1851),
            data_im_in(60) => mul_im_out(1852),
            data_im_in(61) => mul_im_out(1853),
            data_im_in(62) => mul_im_out(1854),
            data_im_in(63) => mul_im_out(1855),
            data_re_out(0) => data_re_out(28),
            data_re_out(1) => data_re_out(60),
            data_re_out(2) => data_re_out(92),
            data_re_out(3) => data_re_out(124),
            data_re_out(4) => data_re_out(156),
            data_re_out(5) => data_re_out(188),
            data_re_out(6) => data_re_out(220),
            data_re_out(7) => data_re_out(252),
            data_re_out(8) => data_re_out(284),
            data_re_out(9) => data_re_out(316),
            data_re_out(10) => data_re_out(348),
            data_re_out(11) => data_re_out(380),
            data_re_out(12) => data_re_out(412),
            data_re_out(13) => data_re_out(444),
            data_re_out(14) => data_re_out(476),
            data_re_out(15) => data_re_out(508),
            data_re_out(16) => data_re_out(540),
            data_re_out(17) => data_re_out(572),
            data_re_out(18) => data_re_out(604),
            data_re_out(19) => data_re_out(636),
            data_re_out(20) => data_re_out(668),
            data_re_out(21) => data_re_out(700),
            data_re_out(22) => data_re_out(732),
            data_re_out(23) => data_re_out(764),
            data_re_out(24) => data_re_out(796),
            data_re_out(25) => data_re_out(828),
            data_re_out(26) => data_re_out(860),
            data_re_out(27) => data_re_out(892),
            data_re_out(28) => data_re_out(924),
            data_re_out(29) => data_re_out(956),
            data_re_out(30) => data_re_out(988),
            data_re_out(31) => data_re_out(1020),
            data_re_out(32) => data_re_out(1052),
            data_re_out(33) => data_re_out(1084),
            data_re_out(34) => data_re_out(1116),
            data_re_out(35) => data_re_out(1148),
            data_re_out(36) => data_re_out(1180),
            data_re_out(37) => data_re_out(1212),
            data_re_out(38) => data_re_out(1244),
            data_re_out(39) => data_re_out(1276),
            data_re_out(40) => data_re_out(1308),
            data_re_out(41) => data_re_out(1340),
            data_re_out(42) => data_re_out(1372),
            data_re_out(43) => data_re_out(1404),
            data_re_out(44) => data_re_out(1436),
            data_re_out(45) => data_re_out(1468),
            data_re_out(46) => data_re_out(1500),
            data_re_out(47) => data_re_out(1532),
            data_re_out(48) => data_re_out(1564),
            data_re_out(49) => data_re_out(1596),
            data_re_out(50) => data_re_out(1628),
            data_re_out(51) => data_re_out(1660),
            data_re_out(52) => data_re_out(1692),
            data_re_out(53) => data_re_out(1724),
            data_re_out(54) => data_re_out(1756),
            data_re_out(55) => data_re_out(1788),
            data_re_out(56) => data_re_out(1820),
            data_re_out(57) => data_re_out(1852),
            data_re_out(58) => data_re_out(1884),
            data_re_out(59) => data_re_out(1916),
            data_re_out(60) => data_re_out(1948),
            data_re_out(61) => data_re_out(1980),
            data_re_out(62) => data_re_out(2012),
            data_re_out(63) => data_re_out(2044),
            data_im_out(0) => data_im_out(28),
            data_im_out(1) => data_im_out(60),
            data_im_out(2) => data_im_out(92),
            data_im_out(3) => data_im_out(124),
            data_im_out(4) => data_im_out(156),
            data_im_out(5) => data_im_out(188),
            data_im_out(6) => data_im_out(220),
            data_im_out(7) => data_im_out(252),
            data_im_out(8) => data_im_out(284),
            data_im_out(9) => data_im_out(316),
            data_im_out(10) => data_im_out(348),
            data_im_out(11) => data_im_out(380),
            data_im_out(12) => data_im_out(412),
            data_im_out(13) => data_im_out(444),
            data_im_out(14) => data_im_out(476),
            data_im_out(15) => data_im_out(508),
            data_im_out(16) => data_im_out(540),
            data_im_out(17) => data_im_out(572),
            data_im_out(18) => data_im_out(604),
            data_im_out(19) => data_im_out(636),
            data_im_out(20) => data_im_out(668),
            data_im_out(21) => data_im_out(700),
            data_im_out(22) => data_im_out(732),
            data_im_out(23) => data_im_out(764),
            data_im_out(24) => data_im_out(796),
            data_im_out(25) => data_im_out(828),
            data_im_out(26) => data_im_out(860),
            data_im_out(27) => data_im_out(892),
            data_im_out(28) => data_im_out(924),
            data_im_out(29) => data_im_out(956),
            data_im_out(30) => data_im_out(988),
            data_im_out(31) => data_im_out(1020),
            data_im_out(32) => data_im_out(1052),
            data_im_out(33) => data_im_out(1084),
            data_im_out(34) => data_im_out(1116),
            data_im_out(35) => data_im_out(1148),
            data_im_out(36) => data_im_out(1180),
            data_im_out(37) => data_im_out(1212),
            data_im_out(38) => data_im_out(1244),
            data_im_out(39) => data_im_out(1276),
            data_im_out(40) => data_im_out(1308),
            data_im_out(41) => data_im_out(1340),
            data_im_out(42) => data_im_out(1372),
            data_im_out(43) => data_im_out(1404),
            data_im_out(44) => data_im_out(1436),
            data_im_out(45) => data_im_out(1468),
            data_im_out(46) => data_im_out(1500),
            data_im_out(47) => data_im_out(1532),
            data_im_out(48) => data_im_out(1564),
            data_im_out(49) => data_im_out(1596),
            data_im_out(50) => data_im_out(1628),
            data_im_out(51) => data_im_out(1660),
            data_im_out(52) => data_im_out(1692),
            data_im_out(53) => data_im_out(1724),
            data_im_out(54) => data_im_out(1756),
            data_im_out(55) => data_im_out(1788),
            data_im_out(56) => data_im_out(1820),
            data_im_out(57) => data_im_out(1852),
            data_im_out(58) => data_im_out(1884),
            data_im_out(59) => data_im_out(1916),
            data_im_out(60) => data_im_out(1948),
            data_im_out(61) => data_im_out(1980),
            data_im_out(62) => data_im_out(2012),
            data_im_out(63) => data_im_out(2044)
        );           

    URFFT_PT64_29 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1856),
            data_re_in(1) => mul_re_out(1857),
            data_re_in(2) => mul_re_out(1858),
            data_re_in(3) => mul_re_out(1859),
            data_re_in(4) => mul_re_out(1860),
            data_re_in(5) => mul_re_out(1861),
            data_re_in(6) => mul_re_out(1862),
            data_re_in(7) => mul_re_out(1863),
            data_re_in(8) => mul_re_out(1864),
            data_re_in(9) => mul_re_out(1865),
            data_re_in(10) => mul_re_out(1866),
            data_re_in(11) => mul_re_out(1867),
            data_re_in(12) => mul_re_out(1868),
            data_re_in(13) => mul_re_out(1869),
            data_re_in(14) => mul_re_out(1870),
            data_re_in(15) => mul_re_out(1871),
            data_re_in(16) => mul_re_out(1872),
            data_re_in(17) => mul_re_out(1873),
            data_re_in(18) => mul_re_out(1874),
            data_re_in(19) => mul_re_out(1875),
            data_re_in(20) => mul_re_out(1876),
            data_re_in(21) => mul_re_out(1877),
            data_re_in(22) => mul_re_out(1878),
            data_re_in(23) => mul_re_out(1879),
            data_re_in(24) => mul_re_out(1880),
            data_re_in(25) => mul_re_out(1881),
            data_re_in(26) => mul_re_out(1882),
            data_re_in(27) => mul_re_out(1883),
            data_re_in(28) => mul_re_out(1884),
            data_re_in(29) => mul_re_out(1885),
            data_re_in(30) => mul_re_out(1886),
            data_re_in(31) => mul_re_out(1887),
            data_re_in(32) => mul_re_out(1888),
            data_re_in(33) => mul_re_out(1889),
            data_re_in(34) => mul_re_out(1890),
            data_re_in(35) => mul_re_out(1891),
            data_re_in(36) => mul_re_out(1892),
            data_re_in(37) => mul_re_out(1893),
            data_re_in(38) => mul_re_out(1894),
            data_re_in(39) => mul_re_out(1895),
            data_re_in(40) => mul_re_out(1896),
            data_re_in(41) => mul_re_out(1897),
            data_re_in(42) => mul_re_out(1898),
            data_re_in(43) => mul_re_out(1899),
            data_re_in(44) => mul_re_out(1900),
            data_re_in(45) => mul_re_out(1901),
            data_re_in(46) => mul_re_out(1902),
            data_re_in(47) => mul_re_out(1903),
            data_re_in(48) => mul_re_out(1904),
            data_re_in(49) => mul_re_out(1905),
            data_re_in(50) => mul_re_out(1906),
            data_re_in(51) => mul_re_out(1907),
            data_re_in(52) => mul_re_out(1908),
            data_re_in(53) => mul_re_out(1909),
            data_re_in(54) => mul_re_out(1910),
            data_re_in(55) => mul_re_out(1911),
            data_re_in(56) => mul_re_out(1912),
            data_re_in(57) => mul_re_out(1913),
            data_re_in(58) => mul_re_out(1914),
            data_re_in(59) => mul_re_out(1915),
            data_re_in(60) => mul_re_out(1916),
            data_re_in(61) => mul_re_out(1917),
            data_re_in(62) => mul_re_out(1918),
            data_re_in(63) => mul_re_out(1919),
            data_im_in(0) => mul_im_out(1856),
            data_im_in(1) => mul_im_out(1857),
            data_im_in(2) => mul_im_out(1858),
            data_im_in(3) => mul_im_out(1859),
            data_im_in(4) => mul_im_out(1860),
            data_im_in(5) => mul_im_out(1861),
            data_im_in(6) => mul_im_out(1862),
            data_im_in(7) => mul_im_out(1863),
            data_im_in(8) => mul_im_out(1864),
            data_im_in(9) => mul_im_out(1865),
            data_im_in(10) => mul_im_out(1866),
            data_im_in(11) => mul_im_out(1867),
            data_im_in(12) => mul_im_out(1868),
            data_im_in(13) => mul_im_out(1869),
            data_im_in(14) => mul_im_out(1870),
            data_im_in(15) => mul_im_out(1871),
            data_im_in(16) => mul_im_out(1872),
            data_im_in(17) => mul_im_out(1873),
            data_im_in(18) => mul_im_out(1874),
            data_im_in(19) => mul_im_out(1875),
            data_im_in(20) => mul_im_out(1876),
            data_im_in(21) => mul_im_out(1877),
            data_im_in(22) => mul_im_out(1878),
            data_im_in(23) => mul_im_out(1879),
            data_im_in(24) => mul_im_out(1880),
            data_im_in(25) => mul_im_out(1881),
            data_im_in(26) => mul_im_out(1882),
            data_im_in(27) => mul_im_out(1883),
            data_im_in(28) => mul_im_out(1884),
            data_im_in(29) => mul_im_out(1885),
            data_im_in(30) => mul_im_out(1886),
            data_im_in(31) => mul_im_out(1887),
            data_im_in(32) => mul_im_out(1888),
            data_im_in(33) => mul_im_out(1889),
            data_im_in(34) => mul_im_out(1890),
            data_im_in(35) => mul_im_out(1891),
            data_im_in(36) => mul_im_out(1892),
            data_im_in(37) => mul_im_out(1893),
            data_im_in(38) => mul_im_out(1894),
            data_im_in(39) => mul_im_out(1895),
            data_im_in(40) => mul_im_out(1896),
            data_im_in(41) => mul_im_out(1897),
            data_im_in(42) => mul_im_out(1898),
            data_im_in(43) => mul_im_out(1899),
            data_im_in(44) => mul_im_out(1900),
            data_im_in(45) => mul_im_out(1901),
            data_im_in(46) => mul_im_out(1902),
            data_im_in(47) => mul_im_out(1903),
            data_im_in(48) => mul_im_out(1904),
            data_im_in(49) => mul_im_out(1905),
            data_im_in(50) => mul_im_out(1906),
            data_im_in(51) => mul_im_out(1907),
            data_im_in(52) => mul_im_out(1908),
            data_im_in(53) => mul_im_out(1909),
            data_im_in(54) => mul_im_out(1910),
            data_im_in(55) => mul_im_out(1911),
            data_im_in(56) => mul_im_out(1912),
            data_im_in(57) => mul_im_out(1913),
            data_im_in(58) => mul_im_out(1914),
            data_im_in(59) => mul_im_out(1915),
            data_im_in(60) => mul_im_out(1916),
            data_im_in(61) => mul_im_out(1917),
            data_im_in(62) => mul_im_out(1918),
            data_im_in(63) => mul_im_out(1919),
            data_re_out(0) => data_re_out(29),
            data_re_out(1) => data_re_out(61),
            data_re_out(2) => data_re_out(93),
            data_re_out(3) => data_re_out(125),
            data_re_out(4) => data_re_out(157),
            data_re_out(5) => data_re_out(189),
            data_re_out(6) => data_re_out(221),
            data_re_out(7) => data_re_out(253),
            data_re_out(8) => data_re_out(285),
            data_re_out(9) => data_re_out(317),
            data_re_out(10) => data_re_out(349),
            data_re_out(11) => data_re_out(381),
            data_re_out(12) => data_re_out(413),
            data_re_out(13) => data_re_out(445),
            data_re_out(14) => data_re_out(477),
            data_re_out(15) => data_re_out(509),
            data_re_out(16) => data_re_out(541),
            data_re_out(17) => data_re_out(573),
            data_re_out(18) => data_re_out(605),
            data_re_out(19) => data_re_out(637),
            data_re_out(20) => data_re_out(669),
            data_re_out(21) => data_re_out(701),
            data_re_out(22) => data_re_out(733),
            data_re_out(23) => data_re_out(765),
            data_re_out(24) => data_re_out(797),
            data_re_out(25) => data_re_out(829),
            data_re_out(26) => data_re_out(861),
            data_re_out(27) => data_re_out(893),
            data_re_out(28) => data_re_out(925),
            data_re_out(29) => data_re_out(957),
            data_re_out(30) => data_re_out(989),
            data_re_out(31) => data_re_out(1021),
            data_re_out(32) => data_re_out(1053),
            data_re_out(33) => data_re_out(1085),
            data_re_out(34) => data_re_out(1117),
            data_re_out(35) => data_re_out(1149),
            data_re_out(36) => data_re_out(1181),
            data_re_out(37) => data_re_out(1213),
            data_re_out(38) => data_re_out(1245),
            data_re_out(39) => data_re_out(1277),
            data_re_out(40) => data_re_out(1309),
            data_re_out(41) => data_re_out(1341),
            data_re_out(42) => data_re_out(1373),
            data_re_out(43) => data_re_out(1405),
            data_re_out(44) => data_re_out(1437),
            data_re_out(45) => data_re_out(1469),
            data_re_out(46) => data_re_out(1501),
            data_re_out(47) => data_re_out(1533),
            data_re_out(48) => data_re_out(1565),
            data_re_out(49) => data_re_out(1597),
            data_re_out(50) => data_re_out(1629),
            data_re_out(51) => data_re_out(1661),
            data_re_out(52) => data_re_out(1693),
            data_re_out(53) => data_re_out(1725),
            data_re_out(54) => data_re_out(1757),
            data_re_out(55) => data_re_out(1789),
            data_re_out(56) => data_re_out(1821),
            data_re_out(57) => data_re_out(1853),
            data_re_out(58) => data_re_out(1885),
            data_re_out(59) => data_re_out(1917),
            data_re_out(60) => data_re_out(1949),
            data_re_out(61) => data_re_out(1981),
            data_re_out(62) => data_re_out(2013),
            data_re_out(63) => data_re_out(2045),
            data_im_out(0) => data_im_out(29),
            data_im_out(1) => data_im_out(61),
            data_im_out(2) => data_im_out(93),
            data_im_out(3) => data_im_out(125),
            data_im_out(4) => data_im_out(157),
            data_im_out(5) => data_im_out(189),
            data_im_out(6) => data_im_out(221),
            data_im_out(7) => data_im_out(253),
            data_im_out(8) => data_im_out(285),
            data_im_out(9) => data_im_out(317),
            data_im_out(10) => data_im_out(349),
            data_im_out(11) => data_im_out(381),
            data_im_out(12) => data_im_out(413),
            data_im_out(13) => data_im_out(445),
            data_im_out(14) => data_im_out(477),
            data_im_out(15) => data_im_out(509),
            data_im_out(16) => data_im_out(541),
            data_im_out(17) => data_im_out(573),
            data_im_out(18) => data_im_out(605),
            data_im_out(19) => data_im_out(637),
            data_im_out(20) => data_im_out(669),
            data_im_out(21) => data_im_out(701),
            data_im_out(22) => data_im_out(733),
            data_im_out(23) => data_im_out(765),
            data_im_out(24) => data_im_out(797),
            data_im_out(25) => data_im_out(829),
            data_im_out(26) => data_im_out(861),
            data_im_out(27) => data_im_out(893),
            data_im_out(28) => data_im_out(925),
            data_im_out(29) => data_im_out(957),
            data_im_out(30) => data_im_out(989),
            data_im_out(31) => data_im_out(1021),
            data_im_out(32) => data_im_out(1053),
            data_im_out(33) => data_im_out(1085),
            data_im_out(34) => data_im_out(1117),
            data_im_out(35) => data_im_out(1149),
            data_im_out(36) => data_im_out(1181),
            data_im_out(37) => data_im_out(1213),
            data_im_out(38) => data_im_out(1245),
            data_im_out(39) => data_im_out(1277),
            data_im_out(40) => data_im_out(1309),
            data_im_out(41) => data_im_out(1341),
            data_im_out(42) => data_im_out(1373),
            data_im_out(43) => data_im_out(1405),
            data_im_out(44) => data_im_out(1437),
            data_im_out(45) => data_im_out(1469),
            data_im_out(46) => data_im_out(1501),
            data_im_out(47) => data_im_out(1533),
            data_im_out(48) => data_im_out(1565),
            data_im_out(49) => data_im_out(1597),
            data_im_out(50) => data_im_out(1629),
            data_im_out(51) => data_im_out(1661),
            data_im_out(52) => data_im_out(1693),
            data_im_out(53) => data_im_out(1725),
            data_im_out(54) => data_im_out(1757),
            data_im_out(55) => data_im_out(1789),
            data_im_out(56) => data_im_out(1821),
            data_im_out(57) => data_im_out(1853),
            data_im_out(58) => data_im_out(1885),
            data_im_out(59) => data_im_out(1917),
            data_im_out(60) => data_im_out(1949),
            data_im_out(61) => data_im_out(1981),
            data_im_out(62) => data_im_out(2013),
            data_im_out(63) => data_im_out(2045)
        );           

    URFFT_PT64_30 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1920),
            data_re_in(1) => mul_re_out(1921),
            data_re_in(2) => mul_re_out(1922),
            data_re_in(3) => mul_re_out(1923),
            data_re_in(4) => mul_re_out(1924),
            data_re_in(5) => mul_re_out(1925),
            data_re_in(6) => mul_re_out(1926),
            data_re_in(7) => mul_re_out(1927),
            data_re_in(8) => mul_re_out(1928),
            data_re_in(9) => mul_re_out(1929),
            data_re_in(10) => mul_re_out(1930),
            data_re_in(11) => mul_re_out(1931),
            data_re_in(12) => mul_re_out(1932),
            data_re_in(13) => mul_re_out(1933),
            data_re_in(14) => mul_re_out(1934),
            data_re_in(15) => mul_re_out(1935),
            data_re_in(16) => mul_re_out(1936),
            data_re_in(17) => mul_re_out(1937),
            data_re_in(18) => mul_re_out(1938),
            data_re_in(19) => mul_re_out(1939),
            data_re_in(20) => mul_re_out(1940),
            data_re_in(21) => mul_re_out(1941),
            data_re_in(22) => mul_re_out(1942),
            data_re_in(23) => mul_re_out(1943),
            data_re_in(24) => mul_re_out(1944),
            data_re_in(25) => mul_re_out(1945),
            data_re_in(26) => mul_re_out(1946),
            data_re_in(27) => mul_re_out(1947),
            data_re_in(28) => mul_re_out(1948),
            data_re_in(29) => mul_re_out(1949),
            data_re_in(30) => mul_re_out(1950),
            data_re_in(31) => mul_re_out(1951),
            data_re_in(32) => mul_re_out(1952),
            data_re_in(33) => mul_re_out(1953),
            data_re_in(34) => mul_re_out(1954),
            data_re_in(35) => mul_re_out(1955),
            data_re_in(36) => mul_re_out(1956),
            data_re_in(37) => mul_re_out(1957),
            data_re_in(38) => mul_re_out(1958),
            data_re_in(39) => mul_re_out(1959),
            data_re_in(40) => mul_re_out(1960),
            data_re_in(41) => mul_re_out(1961),
            data_re_in(42) => mul_re_out(1962),
            data_re_in(43) => mul_re_out(1963),
            data_re_in(44) => mul_re_out(1964),
            data_re_in(45) => mul_re_out(1965),
            data_re_in(46) => mul_re_out(1966),
            data_re_in(47) => mul_re_out(1967),
            data_re_in(48) => mul_re_out(1968),
            data_re_in(49) => mul_re_out(1969),
            data_re_in(50) => mul_re_out(1970),
            data_re_in(51) => mul_re_out(1971),
            data_re_in(52) => mul_re_out(1972),
            data_re_in(53) => mul_re_out(1973),
            data_re_in(54) => mul_re_out(1974),
            data_re_in(55) => mul_re_out(1975),
            data_re_in(56) => mul_re_out(1976),
            data_re_in(57) => mul_re_out(1977),
            data_re_in(58) => mul_re_out(1978),
            data_re_in(59) => mul_re_out(1979),
            data_re_in(60) => mul_re_out(1980),
            data_re_in(61) => mul_re_out(1981),
            data_re_in(62) => mul_re_out(1982),
            data_re_in(63) => mul_re_out(1983),
            data_im_in(0) => mul_im_out(1920),
            data_im_in(1) => mul_im_out(1921),
            data_im_in(2) => mul_im_out(1922),
            data_im_in(3) => mul_im_out(1923),
            data_im_in(4) => mul_im_out(1924),
            data_im_in(5) => mul_im_out(1925),
            data_im_in(6) => mul_im_out(1926),
            data_im_in(7) => mul_im_out(1927),
            data_im_in(8) => mul_im_out(1928),
            data_im_in(9) => mul_im_out(1929),
            data_im_in(10) => mul_im_out(1930),
            data_im_in(11) => mul_im_out(1931),
            data_im_in(12) => mul_im_out(1932),
            data_im_in(13) => mul_im_out(1933),
            data_im_in(14) => mul_im_out(1934),
            data_im_in(15) => mul_im_out(1935),
            data_im_in(16) => mul_im_out(1936),
            data_im_in(17) => mul_im_out(1937),
            data_im_in(18) => mul_im_out(1938),
            data_im_in(19) => mul_im_out(1939),
            data_im_in(20) => mul_im_out(1940),
            data_im_in(21) => mul_im_out(1941),
            data_im_in(22) => mul_im_out(1942),
            data_im_in(23) => mul_im_out(1943),
            data_im_in(24) => mul_im_out(1944),
            data_im_in(25) => mul_im_out(1945),
            data_im_in(26) => mul_im_out(1946),
            data_im_in(27) => mul_im_out(1947),
            data_im_in(28) => mul_im_out(1948),
            data_im_in(29) => mul_im_out(1949),
            data_im_in(30) => mul_im_out(1950),
            data_im_in(31) => mul_im_out(1951),
            data_im_in(32) => mul_im_out(1952),
            data_im_in(33) => mul_im_out(1953),
            data_im_in(34) => mul_im_out(1954),
            data_im_in(35) => mul_im_out(1955),
            data_im_in(36) => mul_im_out(1956),
            data_im_in(37) => mul_im_out(1957),
            data_im_in(38) => mul_im_out(1958),
            data_im_in(39) => mul_im_out(1959),
            data_im_in(40) => mul_im_out(1960),
            data_im_in(41) => mul_im_out(1961),
            data_im_in(42) => mul_im_out(1962),
            data_im_in(43) => mul_im_out(1963),
            data_im_in(44) => mul_im_out(1964),
            data_im_in(45) => mul_im_out(1965),
            data_im_in(46) => mul_im_out(1966),
            data_im_in(47) => mul_im_out(1967),
            data_im_in(48) => mul_im_out(1968),
            data_im_in(49) => mul_im_out(1969),
            data_im_in(50) => mul_im_out(1970),
            data_im_in(51) => mul_im_out(1971),
            data_im_in(52) => mul_im_out(1972),
            data_im_in(53) => mul_im_out(1973),
            data_im_in(54) => mul_im_out(1974),
            data_im_in(55) => mul_im_out(1975),
            data_im_in(56) => mul_im_out(1976),
            data_im_in(57) => mul_im_out(1977),
            data_im_in(58) => mul_im_out(1978),
            data_im_in(59) => mul_im_out(1979),
            data_im_in(60) => mul_im_out(1980),
            data_im_in(61) => mul_im_out(1981),
            data_im_in(62) => mul_im_out(1982),
            data_im_in(63) => mul_im_out(1983),
            data_re_out(0) => data_re_out(30),
            data_re_out(1) => data_re_out(62),
            data_re_out(2) => data_re_out(94),
            data_re_out(3) => data_re_out(126),
            data_re_out(4) => data_re_out(158),
            data_re_out(5) => data_re_out(190),
            data_re_out(6) => data_re_out(222),
            data_re_out(7) => data_re_out(254),
            data_re_out(8) => data_re_out(286),
            data_re_out(9) => data_re_out(318),
            data_re_out(10) => data_re_out(350),
            data_re_out(11) => data_re_out(382),
            data_re_out(12) => data_re_out(414),
            data_re_out(13) => data_re_out(446),
            data_re_out(14) => data_re_out(478),
            data_re_out(15) => data_re_out(510),
            data_re_out(16) => data_re_out(542),
            data_re_out(17) => data_re_out(574),
            data_re_out(18) => data_re_out(606),
            data_re_out(19) => data_re_out(638),
            data_re_out(20) => data_re_out(670),
            data_re_out(21) => data_re_out(702),
            data_re_out(22) => data_re_out(734),
            data_re_out(23) => data_re_out(766),
            data_re_out(24) => data_re_out(798),
            data_re_out(25) => data_re_out(830),
            data_re_out(26) => data_re_out(862),
            data_re_out(27) => data_re_out(894),
            data_re_out(28) => data_re_out(926),
            data_re_out(29) => data_re_out(958),
            data_re_out(30) => data_re_out(990),
            data_re_out(31) => data_re_out(1022),
            data_re_out(32) => data_re_out(1054),
            data_re_out(33) => data_re_out(1086),
            data_re_out(34) => data_re_out(1118),
            data_re_out(35) => data_re_out(1150),
            data_re_out(36) => data_re_out(1182),
            data_re_out(37) => data_re_out(1214),
            data_re_out(38) => data_re_out(1246),
            data_re_out(39) => data_re_out(1278),
            data_re_out(40) => data_re_out(1310),
            data_re_out(41) => data_re_out(1342),
            data_re_out(42) => data_re_out(1374),
            data_re_out(43) => data_re_out(1406),
            data_re_out(44) => data_re_out(1438),
            data_re_out(45) => data_re_out(1470),
            data_re_out(46) => data_re_out(1502),
            data_re_out(47) => data_re_out(1534),
            data_re_out(48) => data_re_out(1566),
            data_re_out(49) => data_re_out(1598),
            data_re_out(50) => data_re_out(1630),
            data_re_out(51) => data_re_out(1662),
            data_re_out(52) => data_re_out(1694),
            data_re_out(53) => data_re_out(1726),
            data_re_out(54) => data_re_out(1758),
            data_re_out(55) => data_re_out(1790),
            data_re_out(56) => data_re_out(1822),
            data_re_out(57) => data_re_out(1854),
            data_re_out(58) => data_re_out(1886),
            data_re_out(59) => data_re_out(1918),
            data_re_out(60) => data_re_out(1950),
            data_re_out(61) => data_re_out(1982),
            data_re_out(62) => data_re_out(2014),
            data_re_out(63) => data_re_out(2046),
            data_im_out(0) => data_im_out(30),
            data_im_out(1) => data_im_out(62),
            data_im_out(2) => data_im_out(94),
            data_im_out(3) => data_im_out(126),
            data_im_out(4) => data_im_out(158),
            data_im_out(5) => data_im_out(190),
            data_im_out(6) => data_im_out(222),
            data_im_out(7) => data_im_out(254),
            data_im_out(8) => data_im_out(286),
            data_im_out(9) => data_im_out(318),
            data_im_out(10) => data_im_out(350),
            data_im_out(11) => data_im_out(382),
            data_im_out(12) => data_im_out(414),
            data_im_out(13) => data_im_out(446),
            data_im_out(14) => data_im_out(478),
            data_im_out(15) => data_im_out(510),
            data_im_out(16) => data_im_out(542),
            data_im_out(17) => data_im_out(574),
            data_im_out(18) => data_im_out(606),
            data_im_out(19) => data_im_out(638),
            data_im_out(20) => data_im_out(670),
            data_im_out(21) => data_im_out(702),
            data_im_out(22) => data_im_out(734),
            data_im_out(23) => data_im_out(766),
            data_im_out(24) => data_im_out(798),
            data_im_out(25) => data_im_out(830),
            data_im_out(26) => data_im_out(862),
            data_im_out(27) => data_im_out(894),
            data_im_out(28) => data_im_out(926),
            data_im_out(29) => data_im_out(958),
            data_im_out(30) => data_im_out(990),
            data_im_out(31) => data_im_out(1022),
            data_im_out(32) => data_im_out(1054),
            data_im_out(33) => data_im_out(1086),
            data_im_out(34) => data_im_out(1118),
            data_im_out(35) => data_im_out(1150),
            data_im_out(36) => data_im_out(1182),
            data_im_out(37) => data_im_out(1214),
            data_im_out(38) => data_im_out(1246),
            data_im_out(39) => data_im_out(1278),
            data_im_out(40) => data_im_out(1310),
            data_im_out(41) => data_im_out(1342),
            data_im_out(42) => data_im_out(1374),
            data_im_out(43) => data_im_out(1406),
            data_im_out(44) => data_im_out(1438),
            data_im_out(45) => data_im_out(1470),
            data_im_out(46) => data_im_out(1502),
            data_im_out(47) => data_im_out(1534),
            data_im_out(48) => data_im_out(1566),
            data_im_out(49) => data_im_out(1598),
            data_im_out(50) => data_im_out(1630),
            data_im_out(51) => data_im_out(1662),
            data_im_out(52) => data_im_out(1694),
            data_im_out(53) => data_im_out(1726),
            data_im_out(54) => data_im_out(1758),
            data_im_out(55) => data_im_out(1790),
            data_im_out(56) => data_im_out(1822),
            data_im_out(57) => data_im_out(1854),
            data_im_out(58) => data_im_out(1886),
            data_im_out(59) => data_im_out(1918),
            data_im_out(60) => data_im_out(1950),
            data_im_out(61) => data_im_out(1982),
            data_im_out(62) => data_im_out(2014),
            data_im_out(63) => data_im_out(2046)
        );           

    URFFT_PT64_31 : fft_pt64
    generic map(
        ctrl_start => (ctrl_start+5) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => (others => '1'),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(1984),
            data_re_in(1) => mul_re_out(1985),
            data_re_in(2) => mul_re_out(1986),
            data_re_in(3) => mul_re_out(1987),
            data_re_in(4) => mul_re_out(1988),
            data_re_in(5) => mul_re_out(1989),
            data_re_in(6) => mul_re_out(1990),
            data_re_in(7) => mul_re_out(1991),
            data_re_in(8) => mul_re_out(1992),
            data_re_in(9) => mul_re_out(1993),
            data_re_in(10) => mul_re_out(1994),
            data_re_in(11) => mul_re_out(1995),
            data_re_in(12) => mul_re_out(1996),
            data_re_in(13) => mul_re_out(1997),
            data_re_in(14) => mul_re_out(1998),
            data_re_in(15) => mul_re_out(1999),
            data_re_in(16) => mul_re_out(2000),
            data_re_in(17) => mul_re_out(2001),
            data_re_in(18) => mul_re_out(2002),
            data_re_in(19) => mul_re_out(2003),
            data_re_in(20) => mul_re_out(2004),
            data_re_in(21) => mul_re_out(2005),
            data_re_in(22) => mul_re_out(2006),
            data_re_in(23) => mul_re_out(2007),
            data_re_in(24) => mul_re_out(2008),
            data_re_in(25) => mul_re_out(2009),
            data_re_in(26) => mul_re_out(2010),
            data_re_in(27) => mul_re_out(2011),
            data_re_in(28) => mul_re_out(2012),
            data_re_in(29) => mul_re_out(2013),
            data_re_in(30) => mul_re_out(2014),
            data_re_in(31) => mul_re_out(2015),
            data_re_in(32) => mul_re_out(2016),
            data_re_in(33) => mul_re_out(2017),
            data_re_in(34) => mul_re_out(2018),
            data_re_in(35) => mul_re_out(2019),
            data_re_in(36) => mul_re_out(2020),
            data_re_in(37) => mul_re_out(2021),
            data_re_in(38) => mul_re_out(2022),
            data_re_in(39) => mul_re_out(2023),
            data_re_in(40) => mul_re_out(2024),
            data_re_in(41) => mul_re_out(2025),
            data_re_in(42) => mul_re_out(2026),
            data_re_in(43) => mul_re_out(2027),
            data_re_in(44) => mul_re_out(2028),
            data_re_in(45) => mul_re_out(2029),
            data_re_in(46) => mul_re_out(2030),
            data_re_in(47) => mul_re_out(2031),
            data_re_in(48) => mul_re_out(2032),
            data_re_in(49) => mul_re_out(2033),
            data_re_in(50) => mul_re_out(2034),
            data_re_in(51) => mul_re_out(2035),
            data_re_in(52) => mul_re_out(2036),
            data_re_in(53) => mul_re_out(2037),
            data_re_in(54) => mul_re_out(2038),
            data_re_in(55) => mul_re_out(2039),
            data_re_in(56) => mul_re_out(2040),
            data_re_in(57) => mul_re_out(2041),
            data_re_in(58) => mul_re_out(2042),
            data_re_in(59) => mul_re_out(2043),
            data_re_in(60) => mul_re_out(2044),
            data_re_in(61) => mul_re_out(2045),
            data_re_in(62) => mul_re_out(2046),
            data_re_in(63) => mul_re_out(2047),
            data_im_in(0) => mul_im_out(1984),
            data_im_in(1) => mul_im_out(1985),
            data_im_in(2) => mul_im_out(1986),
            data_im_in(3) => mul_im_out(1987),
            data_im_in(4) => mul_im_out(1988),
            data_im_in(5) => mul_im_out(1989),
            data_im_in(6) => mul_im_out(1990),
            data_im_in(7) => mul_im_out(1991),
            data_im_in(8) => mul_im_out(1992),
            data_im_in(9) => mul_im_out(1993),
            data_im_in(10) => mul_im_out(1994),
            data_im_in(11) => mul_im_out(1995),
            data_im_in(12) => mul_im_out(1996),
            data_im_in(13) => mul_im_out(1997),
            data_im_in(14) => mul_im_out(1998),
            data_im_in(15) => mul_im_out(1999),
            data_im_in(16) => mul_im_out(2000),
            data_im_in(17) => mul_im_out(2001),
            data_im_in(18) => mul_im_out(2002),
            data_im_in(19) => mul_im_out(2003),
            data_im_in(20) => mul_im_out(2004),
            data_im_in(21) => mul_im_out(2005),
            data_im_in(22) => mul_im_out(2006),
            data_im_in(23) => mul_im_out(2007),
            data_im_in(24) => mul_im_out(2008),
            data_im_in(25) => mul_im_out(2009),
            data_im_in(26) => mul_im_out(2010),
            data_im_in(27) => mul_im_out(2011),
            data_im_in(28) => mul_im_out(2012),
            data_im_in(29) => mul_im_out(2013),
            data_im_in(30) => mul_im_out(2014),
            data_im_in(31) => mul_im_out(2015),
            data_im_in(32) => mul_im_out(2016),
            data_im_in(33) => mul_im_out(2017),
            data_im_in(34) => mul_im_out(2018),
            data_im_in(35) => mul_im_out(2019),
            data_im_in(36) => mul_im_out(2020),
            data_im_in(37) => mul_im_out(2021),
            data_im_in(38) => mul_im_out(2022),
            data_im_in(39) => mul_im_out(2023),
            data_im_in(40) => mul_im_out(2024),
            data_im_in(41) => mul_im_out(2025),
            data_im_in(42) => mul_im_out(2026),
            data_im_in(43) => mul_im_out(2027),
            data_im_in(44) => mul_im_out(2028),
            data_im_in(45) => mul_im_out(2029),
            data_im_in(46) => mul_im_out(2030),
            data_im_in(47) => mul_im_out(2031),
            data_im_in(48) => mul_im_out(2032),
            data_im_in(49) => mul_im_out(2033),
            data_im_in(50) => mul_im_out(2034),
            data_im_in(51) => mul_im_out(2035),
            data_im_in(52) => mul_im_out(2036),
            data_im_in(53) => mul_im_out(2037),
            data_im_in(54) => mul_im_out(2038),
            data_im_in(55) => mul_im_out(2039),
            data_im_in(56) => mul_im_out(2040),
            data_im_in(57) => mul_im_out(2041),
            data_im_in(58) => mul_im_out(2042),
            data_im_in(59) => mul_im_out(2043),
            data_im_in(60) => mul_im_out(2044),
            data_im_in(61) => mul_im_out(2045),
            data_im_in(62) => mul_im_out(2046),
            data_im_in(63) => mul_im_out(2047),
            data_re_out(0) => data_re_out(31),
            data_re_out(1) => data_re_out(63),
            data_re_out(2) => data_re_out(95),
            data_re_out(3) => data_re_out(127),
            data_re_out(4) => data_re_out(159),
            data_re_out(5) => data_re_out(191),
            data_re_out(6) => data_re_out(223),
            data_re_out(7) => data_re_out(255),
            data_re_out(8) => data_re_out(287),
            data_re_out(9) => data_re_out(319),
            data_re_out(10) => data_re_out(351),
            data_re_out(11) => data_re_out(383),
            data_re_out(12) => data_re_out(415),
            data_re_out(13) => data_re_out(447),
            data_re_out(14) => data_re_out(479),
            data_re_out(15) => data_re_out(511),
            data_re_out(16) => data_re_out(543),
            data_re_out(17) => data_re_out(575),
            data_re_out(18) => data_re_out(607),
            data_re_out(19) => data_re_out(639),
            data_re_out(20) => data_re_out(671),
            data_re_out(21) => data_re_out(703),
            data_re_out(22) => data_re_out(735),
            data_re_out(23) => data_re_out(767),
            data_re_out(24) => data_re_out(799),
            data_re_out(25) => data_re_out(831),
            data_re_out(26) => data_re_out(863),
            data_re_out(27) => data_re_out(895),
            data_re_out(28) => data_re_out(927),
            data_re_out(29) => data_re_out(959),
            data_re_out(30) => data_re_out(991),
            data_re_out(31) => data_re_out(1023),
            data_re_out(32) => data_re_out(1055),
            data_re_out(33) => data_re_out(1087),
            data_re_out(34) => data_re_out(1119),
            data_re_out(35) => data_re_out(1151),
            data_re_out(36) => data_re_out(1183),
            data_re_out(37) => data_re_out(1215),
            data_re_out(38) => data_re_out(1247),
            data_re_out(39) => data_re_out(1279),
            data_re_out(40) => data_re_out(1311),
            data_re_out(41) => data_re_out(1343),
            data_re_out(42) => data_re_out(1375),
            data_re_out(43) => data_re_out(1407),
            data_re_out(44) => data_re_out(1439),
            data_re_out(45) => data_re_out(1471),
            data_re_out(46) => data_re_out(1503),
            data_re_out(47) => data_re_out(1535),
            data_re_out(48) => data_re_out(1567),
            data_re_out(49) => data_re_out(1599),
            data_re_out(50) => data_re_out(1631),
            data_re_out(51) => data_re_out(1663),
            data_re_out(52) => data_re_out(1695),
            data_re_out(53) => data_re_out(1727),
            data_re_out(54) => data_re_out(1759),
            data_re_out(55) => data_re_out(1791),
            data_re_out(56) => data_re_out(1823),
            data_re_out(57) => data_re_out(1855),
            data_re_out(58) => data_re_out(1887),
            data_re_out(59) => data_re_out(1919),
            data_re_out(60) => data_re_out(1951),
            data_re_out(61) => data_re_out(1983),
            data_re_out(62) => data_re_out(2015),
            data_re_out(63) => data_re_out(2047),
            data_im_out(0) => data_im_out(31),
            data_im_out(1) => data_im_out(63),
            data_im_out(2) => data_im_out(95),
            data_im_out(3) => data_im_out(127),
            data_im_out(4) => data_im_out(159),
            data_im_out(5) => data_im_out(191),
            data_im_out(6) => data_im_out(223),
            data_im_out(7) => data_im_out(255),
            data_im_out(8) => data_im_out(287),
            data_im_out(9) => data_im_out(319),
            data_im_out(10) => data_im_out(351),
            data_im_out(11) => data_im_out(383),
            data_im_out(12) => data_im_out(415),
            data_im_out(13) => data_im_out(447),
            data_im_out(14) => data_im_out(479),
            data_im_out(15) => data_im_out(511),
            data_im_out(16) => data_im_out(543),
            data_im_out(17) => data_im_out(575),
            data_im_out(18) => data_im_out(607),
            data_im_out(19) => data_im_out(639),
            data_im_out(20) => data_im_out(671),
            data_im_out(21) => data_im_out(703),
            data_im_out(22) => data_im_out(735),
            data_im_out(23) => data_im_out(767),
            data_im_out(24) => data_im_out(799),
            data_im_out(25) => data_im_out(831),
            data_im_out(26) => data_im_out(863),
            data_im_out(27) => data_im_out(895),
            data_im_out(28) => data_im_out(927),
            data_im_out(29) => data_im_out(959),
            data_im_out(30) => data_im_out(991),
            data_im_out(31) => data_im_out(1023),
            data_im_out(32) => data_im_out(1055),
            data_im_out(33) => data_im_out(1087),
            data_im_out(34) => data_im_out(1119),
            data_im_out(35) => data_im_out(1151),
            data_im_out(36) => data_im_out(1183),
            data_im_out(37) => data_im_out(1215),
            data_im_out(38) => data_im_out(1247),
            data_im_out(39) => data_im_out(1279),
            data_im_out(40) => data_im_out(1311),
            data_im_out(41) => data_im_out(1343),
            data_im_out(42) => data_im_out(1375),
            data_im_out(43) => data_im_out(1407),
            data_im_out(44) => data_im_out(1439),
            data_im_out(45) => data_im_out(1471),
            data_im_out(46) => data_im_out(1503),
            data_im_out(47) => data_im_out(1535),
            data_im_out(48) => data_im_out(1567),
            data_im_out(49) => data_im_out(1599),
            data_im_out(50) => data_im_out(1631),
            data_im_out(51) => data_im_out(1663),
            data_im_out(52) => data_im_out(1695),
            data_im_out(53) => data_im_out(1727),
            data_im_out(54) => data_im_out(1759),
            data_im_out(55) => data_im_out(1791),
            data_im_out(56) => data_im_out(1823),
            data_im_out(57) => data_im_out(1855),
            data_im_out(58) => data_im_out(1887),
            data_im_out(59) => data_im_out(1919),
            data_im_out(60) => data_im_out(1951),
            data_im_out(61) => data_im_out(1983),
            data_im_out(62) => data_im_out(2015),
            data_im_out(63) => data_im_out(2047)
        );           


    --- multipliers
 
    UMUL_0 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(0),
            data_im_in => first_stage_im_out(0),
            data_re_out => mul_re_out(0),
            data_im_out => mul_im_out(0)
        );

 
    UMUL_1 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1),
            data_im_in => first_stage_im_out(1),
            data_re_out => mul_re_out(1),
            data_im_out => mul_im_out(1)
        );

 
    UMUL_2 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2),
            data_im_in => first_stage_im_out(2),
            data_re_out => mul_re_out(2),
            data_im_out => mul_im_out(2)
        );

 
    UMUL_3 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(3),
            data_im_in => first_stage_im_out(3),
            data_re_out => mul_re_out(3),
            data_im_out => mul_im_out(3)
        );

 
    UMUL_4 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(4),
            data_im_in => first_stage_im_out(4),
            data_re_out => mul_re_out(4),
            data_im_out => mul_im_out(4)
        );

 
    UMUL_5 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(5),
            data_im_in => first_stage_im_out(5),
            data_re_out => mul_re_out(5),
            data_im_out => mul_im_out(5)
        );

 
    UMUL_6 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(6),
            data_im_in => first_stage_im_out(6),
            data_re_out => mul_re_out(6),
            data_im_out => mul_im_out(6)
        );

 
    UMUL_7 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(7),
            data_im_in => first_stage_im_out(7),
            data_re_out => mul_re_out(7),
            data_im_out => mul_im_out(7)
        );

 
    UMUL_8 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(8),
            data_im_in => first_stage_im_out(8),
            data_re_out => mul_re_out(8),
            data_im_out => mul_im_out(8)
        );

 
    UMUL_9 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(9),
            data_im_in => first_stage_im_out(9),
            data_re_out => mul_re_out(9),
            data_im_out => mul_im_out(9)
        );

 
    UMUL_10 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(10),
            data_im_in => first_stage_im_out(10),
            data_re_out => mul_re_out(10),
            data_im_out => mul_im_out(10)
        );

 
    UMUL_11 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(11),
            data_im_in => first_stage_im_out(11),
            data_re_out => mul_re_out(11),
            data_im_out => mul_im_out(11)
        );

 
    UMUL_12 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(12),
            data_im_in => first_stage_im_out(12),
            data_re_out => mul_re_out(12),
            data_im_out => mul_im_out(12)
        );

 
    UMUL_13 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(13),
            data_im_in => first_stage_im_out(13),
            data_re_out => mul_re_out(13),
            data_im_out => mul_im_out(13)
        );

 
    UMUL_14 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(14),
            data_im_in => first_stage_im_out(14),
            data_re_out => mul_re_out(14),
            data_im_out => mul_im_out(14)
        );

 
    UMUL_15 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(15),
            data_im_in => first_stage_im_out(15),
            data_re_out => mul_re_out(15),
            data_im_out => mul_im_out(15)
        );

 
    UMUL_16 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(16),
            data_im_in => first_stage_im_out(16),
            data_re_out => mul_re_out(16),
            data_im_out => mul_im_out(16)
        );

 
    UMUL_17 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(17),
            data_im_in => first_stage_im_out(17),
            data_re_out => mul_re_out(17),
            data_im_out => mul_im_out(17)
        );

 
    UMUL_18 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(18),
            data_im_in => first_stage_im_out(18),
            data_re_out => mul_re_out(18),
            data_im_out => mul_im_out(18)
        );

 
    UMUL_19 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(19),
            data_im_in => first_stage_im_out(19),
            data_re_out => mul_re_out(19),
            data_im_out => mul_im_out(19)
        );

 
    UMUL_20 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(20),
            data_im_in => first_stage_im_out(20),
            data_re_out => mul_re_out(20),
            data_im_out => mul_im_out(20)
        );

 
    UMUL_21 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(21),
            data_im_in => first_stage_im_out(21),
            data_re_out => mul_re_out(21),
            data_im_out => mul_im_out(21)
        );

 
    UMUL_22 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(22),
            data_im_in => first_stage_im_out(22),
            data_re_out => mul_re_out(22),
            data_im_out => mul_im_out(22)
        );

 
    UMUL_23 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(23),
            data_im_in => first_stage_im_out(23),
            data_re_out => mul_re_out(23),
            data_im_out => mul_im_out(23)
        );

 
    UMUL_24 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(24),
            data_im_in => first_stage_im_out(24),
            data_re_out => mul_re_out(24),
            data_im_out => mul_im_out(24)
        );

 
    UMUL_25 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(25),
            data_im_in => first_stage_im_out(25),
            data_re_out => mul_re_out(25),
            data_im_out => mul_im_out(25)
        );

 
    UMUL_26 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(26),
            data_im_in => first_stage_im_out(26),
            data_re_out => mul_re_out(26),
            data_im_out => mul_im_out(26)
        );

 
    UMUL_27 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(27),
            data_im_in => first_stage_im_out(27),
            data_re_out => mul_re_out(27),
            data_im_out => mul_im_out(27)
        );

 
    UMUL_28 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(28),
            data_im_in => first_stage_im_out(28),
            data_re_out => mul_re_out(28),
            data_im_out => mul_im_out(28)
        );

 
    UMUL_29 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(29),
            data_im_in => first_stage_im_out(29),
            data_re_out => mul_re_out(29),
            data_im_out => mul_im_out(29)
        );

 
    UMUL_30 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(30),
            data_im_in => first_stage_im_out(30),
            data_re_out => mul_re_out(30),
            data_im_out => mul_im_out(30)
        );

 
    UMUL_31 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(31),
            data_im_in => first_stage_im_out(31),
            data_re_out => mul_re_out(31),
            data_im_out => mul_im_out(31)
        );

 
    UMUL_32 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(32),
            data_im_in => first_stage_im_out(32),
            data_re_out => mul_re_out(32),
            data_im_out => mul_im_out(32)
        );

 
    UMUL_33 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(33),
            data_im_in => first_stage_im_out(33),
            data_re_out => mul_re_out(33),
            data_im_out => mul_im_out(33)
        );

 
    UMUL_34 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(34),
            data_im_in => first_stage_im_out(34),
            data_re_out => mul_re_out(34),
            data_im_out => mul_im_out(34)
        );

 
    UMUL_35 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(35),
            data_im_in => first_stage_im_out(35),
            data_re_out => mul_re_out(35),
            data_im_out => mul_im_out(35)
        );

 
    UMUL_36 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(36),
            data_im_in => first_stage_im_out(36),
            data_re_out => mul_re_out(36),
            data_im_out => mul_im_out(36)
        );

 
    UMUL_37 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(37),
            data_im_in => first_stage_im_out(37),
            data_re_out => mul_re_out(37),
            data_im_out => mul_im_out(37)
        );

 
    UMUL_38 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(38),
            data_im_in => first_stage_im_out(38),
            data_re_out => mul_re_out(38),
            data_im_out => mul_im_out(38)
        );

 
    UMUL_39 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(39),
            data_im_in => first_stage_im_out(39),
            data_re_out => mul_re_out(39),
            data_im_out => mul_im_out(39)
        );

 
    UMUL_40 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(40),
            data_im_in => first_stage_im_out(40),
            data_re_out => mul_re_out(40),
            data_im_out => mul_im_out(40)
        );

 
    UMUL_41 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(41),
            data_im_in => first_stage_im_out(41),
            data_re_out => mul_re_out(41),
            data_im_out => mul_im_out(41)
        );

 
    UMUL_42 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(42),
            data_im_in => first_stage_im_out(42),
            data_re_out => mul_re_out(42),
            data_im_out => mul_im_out(42)
        );

 
    UMUL_43 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(43),
            data_im_in => first_stage_im_out(43),
            data_re_out => mul_re_out(43),
            data_im_out => mul_im_out(43)
        );

 
    UMUL_44 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(44),
            data_im_in => first_stage_im_out(44),
            data_re_out => mul_re_out(44),
            data_im_out => mul_im_out(44)
        );

 
    UMUL_45 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(45),
            data_im_in => first_stage_im_out(45),
            data_re_out => mul_re_out(45),
            data_im_out => mul_im_out(45)
        );

 
    UMUL_46 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(46),
            data_im_in => first_stage_im_out(46),
            data_re_out => mul_re_out(46),
            data_im_out => mul_im_out(46)
        );

 
    UMUL_47 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(47),
            data_im_in => first_stage_im_out(47),
            data_re_out => mul_re_out(47),
            data_im_out => mul_im_out(47)
        );

 
    UMUL_48 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(48),
            data_im_in => first_stage_im_out(48),
            data_re_out => mul_re_out(48),
            data_im_out => mul_im_out(48)
        );

 
    UMUL_49 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(49),
            data_im_in => first_stage_im_out(49),
            data_re_out => mul_re_out(49),
            data_im_out => mul_im_out(49)
        );

 
    UMUL_50 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(50),
            data_im_in => first_stage_im_out(50),
            data_re_out => mul_re_out(50),
            data_im_out => mul_im_out(50)
        );

 
    UMUL_51 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(51),
            data_im_in => first_stage_im_out(51),
            data_re_out => mul_re_out(51),
            data_im_out => mul_im_out(51)
        );

 
    UMUL_52 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(52),
            data_im_in => first_stage_im_out(52),
            data_re_out => mul_re_out(52),
            data_im_out => mul_im_out(52)
        );

 
    UMUL_53 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(53),
            data_im_in => first_stage_im_out(53),
            data_re_out => mul_re_out(53),
            data_im_out => mul_im_out(53)
        );

 
    UMUL_54 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(54),
            data_im_in => first_stage_im_out(54),
            data_re_out => mul_re_out(54),
            data_im_out => mul_im_out(54)
        );

 
    UMUL_55 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(55),
            data_im_in => first_stage_im_out(55),
            data_re_out => mul_re_out(55),
            data_im_out => mul_im_out(55)
        );

 
    UMUL_56 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(56),
            data_im_in => first_stage_im_out(56),
            data_re_out => mul_re_out(56),
            data_im_out => mul_im_out(56)
        );

 
    UMUL_57 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(57),
            data_im_in => first_stage_im_out(57),
            data_re_out => mul_re_out(57),
            data_im_out => mul_im_out(57)
        );

 
    UMUL_58 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(58),
            data_im_in => first_stage_im_out(58),
            data_re_out => mul_re_out(58),
            data_im_out => mul_im_out(58)
        );

 
    UMUL_59 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(59),
            data_im_in => first_stage_im_out(59),
            data_re_out => mul_re_out(59),
            data_im_out => mul_im_out(59)
        );

 
    UMUL_60 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(60),
            data_im_in => first_stage_im_out(60),
            data_re_out => mul_re_out(60),
            data_im_out => mul_im_out(60)
        );

 
    UMUL_61 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(61),
            data_im_in => first_stage_im_out(61),
            data_re_out => mul_re_out(61),
            data_im_out => mul_im_out(61)
        );

 
    UMUL_62 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(62),
            data_im_in => first_stage_im_out(62),
            data_re_out => mul_re_out(62),
            data_im_out => mul_im_out(62)
        );

 
    UMUL_63 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(63),
            data_im_in => first_stage_im_out(63),
            data_re_out => mul_re_out(63),
            data_im_out => mul_im_out(63)
        );

 
    UMUL_64 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(64),
            data_im_in => first_stage_im_out(64),
            data_re_out => mul_re_out(64),
            data_im_out => mul_im_out(64)
        );

 
    UMUL_65 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(65),
            data_im_in => first_stage_im_out(65),
            re_multiplicator => "0100000000000000", --- 1.0 + j-0.0030517578125
            im_multiplicator => "1111111111001110",
            data_re_out => mul_re_out(65),
            data_im_out => mul_im_out(65)
        );

 
    UMUL_66 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(66),
            data_im_in => first_stage_im_out(66),
            re_multiplicator => "0100000000000000", --- 1.0 + j-0.00616455078125
            im_multiplicator => "1111111110011011",
            data_re_out => mul_re_out(66),
            data_im_out => mul_im_out(66)
        );

 
    UMUL_67 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(67),
            data_im_in => first_stage_im_out(67),
            re_multiplicator => "0011111111111111", --- 0.999938964844 + j-0.00921630859375
            im_multiplicator => "1111111101101001",
            data_re_out => mul_re_out(67),
            data_im_out => mul_im_out(67)
        );

 
    UMUL_68 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(68),
            data_im_in => first_stage_im_out(68),
            re_multiplicator => "0011111111111111", --- 0.999938964844 + j-0.0122680664062
            im_multiplicator => "1111111100110111",
            data_re_out => mul_re_out(68),
            data_im_out => mul_im_out(68)
        );

 
    UMUL_69 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(69),
            data_im_in => first_stage_im_out(69),
            re_multiplicator => "0011111111111110", --- 0.999877929688 + j-0.0153198242188
            im_multiplicator => "1111111100000101",
            data_re_out => mul_re_out(69),
            data_im_out => mul_im_out(69)
        );

 
    UMUL_70 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(70),
            data_im_in => first_stage_im_out(70),
            re_multiplicator => "0011111111111101", --- 0.999816894531 + j-0.0184326171875
            im_multiplicator => "1111111011010010",
            data_re_out => mul_re_out(70),
            data_im_out => mul_im_out(70)
        );

 
    UMUL_71 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(71),
            data_im_in => first_stage_im_out(71),
            re_multiplicator => "0011111111111100", --- 0.999755859375 + j-0.021484375
            im_multiplicator => "1111111010100000",
            data_re_out => mul_re_out(71),
            data_im_out => mul_im_out(71)
        );

 
    UMUL_72 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(72),
            data_im_in => first_stage_im_out(72),
            re_multiplicator => "0011111111111011", --- 0.999694824219 + j-0.0245361328125
            im_multiplicator => "1111111001101110",
            data_re_out => mul_re_out(72),
            data_im_out => mul_im_out(72)
        );

 
    UMUL_73 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(73),
            data_im_in => first_stage_im_out(73),
            re_multiplicator => "0011111111111010", --- 0.999633789062 + j-0.027587890625
            im_multiplicator => "1111111000111100",
            data_re_out => mul_re_out(73),
            data_im_out => mul_im_out(73)
        );

 
    UMUL_74 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(74),
            data_im_in => first_stage_im_out(74),
            re_multiplicator => "0011111111111000", --- 0.99951171875 + j-0.0307006835938
            im_multiplicator => "1111111000001001",
            data_re_out => mul_re_out(74),
            data_im_out => mul_im_out(74)
        );

 
    UMUL_75 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(75),
            data_im_in => first_stage_im_out(75),
            re_multiplicator => "0011111111110111", --- 0.999450683594 + j-0.0337524414062
            im_multiplicator => "1111110111010111",
            data_re_out => mul_re_out(75),
            data_im_out => mul_im_out(75)
        );

 
    UMUL_76 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(76),
            data_im_in => first_stage_im_out(76),
            re_multiplicator => "0011111111110101", --- 0.999328613281 + j-0.0368041992188
            im_multiplicator => "1111110110100101",
            data_re_out => mul_re_out(76),
            data_im_out => mul_im_out(76)
        );

 
    UMUL_77 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(77),
            data_im_in => first_stage_im_out(77),
            re_multiplicator => "0011111111110011", --- 0.999206542969 + j-0.0398559570312
            im_multiplicator => "1111110101110011",
            data_re_out => mul_re_out(77),
            data_im_out => mul_im_out(77)
        );

 
    UMUL_78 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(78),
            data_im_in => first_stage_im_out(78),
            re_multiplicator => "0011111111110001", --- 0.999084472656 + j-0.04296875
            im_multiplicator => "1111110101000000",
            data_re_out => mul_re_out(78),
            data_im_out => mul_im_out(78)
        );

 
    UMUL_79 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(79),
            data_im_in => first_stage_im_out(79),
            re_multiplicator => "0011111111101111", --- 0.998962402344 + j-0.0460205078125
            im_multiplicator => "1111110100001110",
            data_re_out => mul_re_out(79),
            data_im_out => mul_im_out(79)
        );

 
    UMUL_80 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(80),
            data_im_in => first_stage_im_out(80),
            re_multiplicator => "0011111111101100", --- 0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(80),
            data_im_out => mul_im_out(80)
        );

 
    UMUL_81 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(81),
            data_im_in => first_stage_im_out(81),
            re_multiplicator => "0011111111101010", --- 0.998657226562 + j-0.0521240234375
            im_multiplicator => "1111110010101010",
            data_re_out => mul_re_out(81),
            data_im_out => mul_im_out(81)
        );

 
    UMUL_82 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(82),
            data_im_in => first_stage_im_out(82),
            re_multiplicator => "0011111111100111", --- 0.998474121094 + j-0.05517578125
            im_multiplicator => "1111110001111000",
            data_re_out => mul_re_out(82),
            data_im_out => mul_im_out(82)
        );

 
    UMUL_83 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(83),
            data_im_in => first_stage_im_out(83),
            re_multiplicator => "0011111111100100", --- 0.998291015625 + j-0.0582885742188
            im_multiplicator => "1111110001000101",
            data_re_out => mul_re_out(83),
            data_im_out => mul_im_out(83)
        );

 
    UMUL_84 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(84),
            data_im_in => first_stage_im_out(84),
            re_multiplicator => "0011111111100001", --- 0.998107910156 + j-0.0613403320312
            im_multiplicator => "1111110000010011",
            data_re_out => mul_re_out(84),
            data_im_out => mul_im_out(84)
        );

 
    UMUL_85 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(85),
            data_im_in => first_stage_im_out(85),
            re_multiplicator => "0011111111011110", --- 0.997924804688 + j-0.0643920898438
            im_multiplicator => "1111101111100001",
            data_re_out => mul_re_out(85),
            data_im_out => mul_im_out(85)
        );

 
    UMUL_86 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(86),
            data_im_in => first_stage_im_out(86),
            re_multiplicator => "0011111111011011", --- 0.997741699219 + j-0.0674438476562
            im_multiplicator => "1111101110101111",
            data_re_out => mul_re_out(86),
            data_im_out => mul_im_out(86)
        );

 
    UMUL_87 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(87),
            data_im_in => first_stage_im_out(87),
            re_multiplicator => "0011111111010111", --- 0.997497558594 + j-0.0704956054688
            im_multiplicator => "1111101101111101",
            data_re_out => mul_re_out(87),
            data_im_out => mul_im_out(87)
        );

 
    UMUL_88 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(88),
            data_im_in => first_stage_im_out(88),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(88),
            data_im_out => mul_im_out(88)
        );

 
    UMUL_89 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(89),
            data_im_in => first_stage_im_out(89),
            re_multiplicator => "0011111111010000", --- 0.9970703125 + j-0.0765991210938
            im_multiplicator => "1111101100011001",
            data_re_out => mul_re_out(89),
            data_im_out => mul_im_out(89)
        );

 
    UMUL_90 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(90),
            data_im_in => first_stage_im_out(90),
            re_multiplicator => "0011111111001100", --- 0.996826171875 + j-0.0797119140625
            im_multiplicator => "1111101011100110",
            data_re_out => mul_re_out(90),
            data_im_out => mul_im_out(90)
        );

 
    UMUL_91 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(91),
            data_im_in => first_stage_im_out(91),
            re_multiplicator => "0011111111001000", --- 0.99658203125 + j-0.082763671875
            im_multiplicator => "1111101010110100",
            data_re_out => mul_re_out(91),
            data_im_out => mul_im_out(91)
        );

 
    UMUL_92 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(92),
            data_im_in => first_stage_im_out(92),
            re_multiplicator => "0011111111000100", --- 0.996337890625 + j-0.0858154296875
            im_multiplicator => "1111101010000010",
            data_re_out => mul_re_out(92),
            data_im_out => mul_im_out(92)
        );

 
    UMUL_93 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(93),
            data_im_in => first_stage_im_out(93),
            re_multiplicator => "0011111110111111", --- 0.996032714844 + j-0.0888671875
            im_multiplicator => "1111101001010000",
            data_re_out => mul_re_out(93),
            data_im_out => mul_im_out(93)
        );

 
    UMUL_94 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(94),
            data_im_in => first_stage_im_out(94),
            re_multiplicator => "0011111110111011", --- 0.995788574219 + j-0.0919189453125
            im_multiplicator => "1111101000011110",
            data_re_out => mul_re_out(94),
            data_im_out => mul_im_out(94)
        );

 
    UMUL_95 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(95),
            data_im_in => first_stage_im_out(95),
            re_multiplicator => "0011111110110110", --- 0.995483398438 + j-0.094970703125
            im_multiplicator => "1111100111101100",
            data_re_out => mul_re_out(95),
            data_im_out => mul_im_out(95)
        );

 
    UMUL_96 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(96),
            data_im_in => first_stage_im_out(96),
            re_multiplicator => "0011111110110001", --- 0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(96),
            data_im_out => mul_im_out(96)
        );

 
    UMUL_97 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(97),
            data_im_in => first_stage_im_out(97),
            re_multiplicator => "0011111110101100", --- 0.994873046875 + j-0.10107421875
            im_multiplicator => "1111100110001000",
            data_re_out => mul_re_out(97),
            data_im_out => mul_im_out(97)
        );

 
    UMUL_98 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(98),
            data_im_in => first_stage_im_out(98),
            re_multiplicator => "0011111110100111", --- 0.994567871094 + j-0.104125976562
            im_multiplicator => "1111100101010110",
            data_re_out => mul_re_out(98),
            data_im_out => mul_im_out(98)
        );

 
    UMUL_99 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(99),
            data_im_in => first_stage_im_out(99),
            re_multiplicator => "0011111110100010", --- 0.994262695312 + j-0.107177734375
            im_multiplicator => "1111100100100100",
            data_re_out => mul_re_out(99),
            data_im_out => mul_im_out(99)
        );

 
    UMUL_100 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(100),
            data_im_in => first_stage_im_out(100),
            re_multiplicator => "0011111110011100", --- 0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(100),
            data_im_out => mul_im_out(100)
        );

 
    UMUL_101 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(101),
            data_im_in => first_stage_im_out(101),
            re_multiplicator => "0011111110010111", --- 0.993591308594 + j-0.11328125
            im_multiplicator => "1111100011000000",
            data_re_out => mul_re_out(101),
            data_im_out => mul_im_out(101)
        );

 
    UMUL_102 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(102),
            data_im_in => first_stage_im_out(102),
            re_multiplicator => "0011111110010001", --- 0.993225097656 + j-0.116333007812
            im_multiplicator => "1111100010001110",
            data_re_out => mul_re_out(102),
            data_im_out => mul_im_out(102)
        );

 
    UMUL_103 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(103),
            data_im_in => first_stage_im_out(103),
            re_multiplicator => "0011111110001011", --- 0.992858886719 + j-0.119384765625
            im_multiplicator => "1111100001011100",
            data_re_out => mul_re_out(103),
            data_im_out => mul_im_out(103)
        );

 
    UMUL_104 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(104),
            data_im_in => first_stage_im_out(104),
            re_multiplicator => "0011111110000101", --- 0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(104),
            data_im_out => mul_im_out(104)
        );

 
    UMUL_105 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(105),
            data_im_in => first_stage_im_out(105),
            re_multiplicator => "0011111101111111", --- 0.992126464844 + j-0.125427246094
            im_multiplicator => "1111011111111001",
            data_re_out => mul_re_out(105),
            data_im_out => mul_im_out(105)
        );

 
    UMUL_106 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(106),
            data_im_in => first_stage_im_out(106),
            re_multiplicator => "0011111101111000", --- 0.99169921875 + j-0.128479003906
            im_multiplicator => "1111011111000111",
            data_re_out => mul_re_out(106),
            data_im_out => mul_im_out(106)
        );

 
    UMUL_107 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(107),
            data_im_in => first_stage_im_out(107),
            re_multiplicator => "0011111101110010", --- 0.991333007812 + j-0.131530761719
            im_multiplicator => "1111011110010101",
            data_re_out => mul_re_out(107),
            data_im_out => mul_im_out(107)
        );

 
    UMUL_108 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(108),
            data_im_in => first_stage_im_out(108),
            re_multiplicator => "0011111101101011", --- 0.990905761719 + j-0.134582519531
            im_multiplicator => "1111011101100011",
            data_re_out => mul_re_out(108),
            data_im_out => mul_im_out(108)
        );

 
    UMUL_109 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(109),
            data_im_in => first_stage_im_out(109),
            re_multiplicator => "0011111101100100", --- 0.990478515625 + j-0.137634277344
            im_multiplicator => "1111011100110001",
            data_re_out => mul_re_out(109),
            data_im_out => mul_im_out(109)
        );

 
    UMUL_110 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(110),
            data_im_in => first_stage_im_out(110),
            re_multiplicator => "0011111101011101", --- 0.990051269531 + j-0.140686035156
            im_multiplicator => "1111011011111111",
            data_re_out => mul_re_out(110),
            data_im_out => mul_im_out(110)
        );

 
    UMUL_111 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(111),
            data_im_in => first_stage_im_out(111),
            re_multiplicator => "0011111101010110", --- 0.989624023438 + j-0.143676757812
            im_multiplicator => "1111011011001110",
            data_re_out => mul_re_out(111),
            data_im_out => mul_im_out(111)
        );

 
    UMUL_112 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(112),
            data_im_in => first_stage_im_out(112),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(112),
            data_im_out => mul_im_out(112)
        );

 
    UMUL_113 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(113),
            data_im_in => first_stage_im_out(113),
            re_multiplicator => "0011111101000111", --- 0.988708496094 + j-0.149780273438
            im_multiplicator => "1111011001101010",
            data_re_out => mul_re_out(113),
            data_im_out => mul_im_out(113)
        );

 
    UMUL_114 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(114),
            data_im_in => first_stage_im_out(114),
            re_multiplicator => "0011111101000000", --- 0.98828125 + j-0.152770996094
            im_multiplicator => "1111011000111001",
            data_re_out => mul_re_out(114),
            data_im_out => mul_im_out(114)
        );

 
    UMUL_115 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(115),
            data_im_in => first_stage_im_out(115),
            re_multiplicator => "0011111100111000", --- 0.98779296875 + j-0.155822753906
            im_multiplicator => "1111011000000111",
            data_re_out => mul_re_out(115),
            data_im_out => mul_im_out(115)
        );

 
    UMUL_116 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(116),
            data_im_in => first_stage_im_out(116),
            re_multiplicator => "0011111100110000", --- 0.9873046875 + j-0.158874511719
            im_multiplicator => "1111010111010101",
            data_re_out => mul_re_out(116),
            data_im_out => mul_im_out(116)
        );

 
    UMUL_117 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(117),
            data_im_in => first_stage_im_out(117),
            re_multiplicator => "0011111100101000", --- 0.98681640625 + j-0.161865234375
            im_multiplicator => "1111010110100100",
            data_re_out => mul_re_out(117),
            data_im_out => mul_im_out(117)
        );

 
    UMUL_118 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(118),
            data_im_in => first_stage_im_out(118),
            re_multiplicator => "0011111100100000", --- 0.986328125 + j-0.164916992188
            im_multiplicator => "1111010101110010",
            data_re_out => mul_re_out(118),
            data_im_out => mul_im_out(118)
        );

 
    UMUL_119 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(119),
            data_im_in => first_stage_im_out(119),
            re_multiplicator => "0011111100010111", --- 0.985778808594 + j-0.16796875
            im_multiplicator => "1111010101000000",
            data_re_out => mul_re_out(119),
            data_im_out => mul_im_out(119)
        );

 
    UMUL_120 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(120),
            data_im_in => first_stage_im_out(120),
            re_multiplicator => "0011111100001111", --- 0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(120),
            data_im_out => mul_im_out(120)
        );

 
    UMUL_121 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(121),
            data_im_in => first_stage_im_out(121),
            re_multiplicator => "0011111100000110", --- 0.984741210938 + j-0.174011230469
            im_multiplicator => "1111010011011101",
            data_re_out => mul_re_out(121),
            data_im_out => mul_im_out(121)
        );

 
    UMUL_122 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(122),
            data_im_in => first_stage_im_out(122),
            re_multiplicator => "0011111011111101", --- 0.984191894531 + j-0.177001953125
            im_multiplicator => "1111010010101100",
            data_re_out => mul_re_out(122),
            data_im_out => mul_im_out(122)
        );

 
    UMUL_123 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(123),
            data_im_in => first_stage_im_out(123),
            re_multiplicator => "0011111011110100", --- 0.983642578125 + j-0.179992675781
            im_multiplicator => "1111010001111011",
            data_re_out => mul_re_out(123),
            data_im_out => mul_im_out(123)
        );

 
    UMUL_124 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(124),
            data_im_in => first_stage_im_out(124),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(124),
            data_im_out => mul_im_out(124)
        );

 
    UMUL_125 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(125),
            data_im_in => first_stage_im_out(125),
            re_multiplicator => "0011111011100010", --- 0.982543945312 + j-0.18603515625
            im_multiplicator => "1111010000011000",
            data_re_out => mul_re_out(125),
            data_im_out => mul_im_out(125)
        );

 
    UMUL_126 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(126),
            data_im_in => first_stage_im_out(126),
            re_multiplicator => "0011111011011000", --- 0.98193359375 + j-0.189086914062
            im_multiplicator => "1111001111100110",
            data_re_out => mul_re_out(126),
            data_im_out => mul_im_out(126)
        );

 
    UMUL_127 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(127),
            data_im_in => first_stage_im_out(127),
            re_multiplicator => "0011111011001111", --- 0.981384277344 + j-0.192077636719
            im_multiplicator => "1111001110110101",
            data_re_out => mul_re_out(127),
            data_im_out => mul_im_out(127)
        );

 
    UMUL_128 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(128),
            data_im_in => first_stage_im_out(128),
            data_re_out => mul_re_out(128),
            data_im_out => mul_im_out(128)
        );

 
    UMUL_129 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(129),
            data_im_in => first_stage_im_out(129),
            re_multiplicator => "0100000000000000", --- 1.0 + j-0.00616455078125
            im_multiplicator => "1111111110011011",
            data_re_out => mul_re_out(129),
            data_im_out => mul_im_out(129)
        );

 
    UMUL_130 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(130),
            data_im_in => first_stage_im_out(130),
            re_multiplicator => "0011111111111111", --- 0.999938964844 + j-0.0122680664062
            im_multiplicator => "1111111100110111",
            data_re_out => mul_re_out(130),
            data_im_out => mul_im_out(130)
        );

 
    UMUL_131 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(131),
            data_im_in => first_stage_im_out(131),
            re_multiplicator => "0011111111111101", --- 0.999816894531 + j-0.0184326171875
            im_multiplicator => "1111111011010010",
            data_re_out => mul_re_out(131),
            data_im_out => mul_im_out(131)
        );

 
    UMUL_132 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(132),
            data_im_in => first_stage_im_out(132),
            re_multiplicator => "0011111111111011", --- 0.999694824219 + j-0.0245361328125
            im_multiplicator => "1111111001101110",
            data_re_out => mul_re_out(132),
            data_im_out => mul_im_out(132)
        );

 
    UMUL_133 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(133),
            data_im_in => first_stage_im_out(133),
            re_multiplicator => "0011111111111000", --- 0.99951171875 + j-0.0307006835938
            im_multiplicator => "1111111000001001",
            data_re_out => mul_re_out(133),
            data_im_out => mul_im_out(133)
        );

 
    UMUL_134 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(134),
            data_im_in => first_stage_im_out(134),
            re_multiplicator => "0011111111110101", --- 0.999328613281 + j-0.0368041992188
            im_multiplicator => "1111110110100101",
            data_re_out => mul_re_out(134),
            data_im_out => mul_im_out(134)
        );

 
    UMUL_135 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(135),
            data_im_in => first_stage_im_out(135),
            re_multiplicator => "0011111111110001", --- 0.999084472656 + j-0.04296875
            im_multiplicator => "1111110101000000",
            data_re_out => mul_re_out(135),
            data_im_out => mul_im_out(135)
        );

 
    UMUL_136 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(136),
            data_im_in => first_stage_im_out(136),
            re_multiplicator => "0011111111101100", --- 0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(136),
            data_im_out => mul_im_out(136)
        );

 
    UMUL_137 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(137),
            data_im_in => first_stage_im_out(137),
            re_multiplicator => "0011111111100111", --- 0.998474121094 + j-0.05517578125
            im_multiplicator => "1111110001111000",
            data_re_out => mul_re_out(137),
            data_im_out => mul_im_out(137)
        );

 
    UMUL_138 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(138),
            data_im_in => first_stage_im_out(138),
            re_multiplicator => "0011111111100001", --- 0.998107910156 + j-0.0613403320312
            im_multiplicator => "1111110000010011",
            data_re_out => mul_re_out(138),
            data_im_out => mul_im_out(138)
        );

 
    UMUL_139 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(139),
            data_im_in => first_stage_im_out(139),
            re_multiplicator => "0011111111011011", --- 0.997741699219 + j-0.0674438476562
            im_multiplicator => "1111101110101111",
            data_re_out => mul_re_out(139),
            data_im_out => mul_im_out(139)
        );

 
    UMUL_140 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(140),
            data_im_in => first_stage_im_out(140),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(140),
            data_im_out => mul_im_out(140)
        );

 
    UMUL_141 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(141),
            data_im_in => first_stage_im_out(141),
            re_multiplicator => "0011111111001100", --- 0.996826171875 + j-0.0797119140625
            im_multiplicator => "1111101011100110",
            data_re_out => mul_re_out(141),
            data_im_out => mul_im_out(141)
        );

 
    UMUL_142 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(142),
            data_im_in => first_stage_im_out(142),
            re_multiplicator => "0011111111000100", --- 0.996337890625 + j-0.0858154296875
            im_multiplicator => "1111101010000010",
            data_re_out => mul_re_out(142),
            data_im_out => mul_im_out(142)
        );

 
    UMUL_143 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(143),
            data_im_in => first_stage_im_out(143),
            re_multiplicator => "0011111110111011", --- 0.995788574219 + j-0.0919189453125
            im_multiplicator => "1111101000011110",
            data_re_out => mul_re_out(143),
            data_im_out => mul_im_out(143)
        );

 
    UMUL_144 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(144),
            data_im_in => first_stage_im_out(144),
            re_multiplicator => "0011111110110001", --- 0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(144),
            data_im_out => mul_im_out(144)
        );

 
    UMUL_145 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(145),
            data_im_in => first_stage_im_out(145),
            re_multiplicator => "0011111110100111", --- 0.994567871094 + j-0.104125976562
            im_multiplicator => "1111100101010110",
            data_re_out => mul_re_out(145),
            data_im_out => mul_im_out(145)
        );

 
    UMUL_146 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(146),
            data_im_in => first_stage_im_out(146),
            re_multiplicator => "0011111110011100", --- 0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(146),
            data_im_out => mul_im_out(146)
        );

 
    UMUL_147 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(147),
            data_im_in => first_stage_im_out(147),
            re_multiplicator => "0011111110010001", --- 0.993225097656 + j-0.116333007812
            im_multiplicator => "1111100010001110",
            data_re_out => mul_re_out(147),
            data_im_out => mul_im_out(147)
        );

 
    UMUL_148 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(148),
            data_im_in => first_stage_im_out(148),
            re_multiplicator => "0011111110000101", --- 0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(148),
            data_im_out => mul_im_out(148)
        );

 
    UMUL_149 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(149),
            data_im_in => first_stage_im_out(149),
            re_multiplicator => "0011111101111000", --- 0.99169921875 + j-0.128479003906
            im_multiplicator => "1111011111000111",
            data_re_out => mul_re_out(149),
            data_im_out => mul_im_out(149)
        );

 
    UMUL_150 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(150),
            data_im_in => first_stage_im_out(150),
            re_multiplicator => "0011111101101011", --- 0.990905761719 + j-0.134582519531
            im_multiplicator => "1111011101100011",
            data_re_out => mul_re_out(150),
            data_im_out => mul_im_out(150)
        );

 
    UMUL_151 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(151),
            data_im_in => first_stage_im_out(151),
            re_multiplicator => "0011111101011101", --- 0.990051269531 + j-0.140686035156
            im_multiplicator => "1111011011111111",
            data_re_out => mul_re_out(151),
            data_im_out => mul_im_out(151)
        );

 
    UMUL_152 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(152),
            data_im_in => first_stage_im_out(152),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(152),
            data_im_out => mul_im_out(152)
        );

 
    UMUL_153 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(153),
            data_im_in => first_stage_im_out(153),
            re_multiplicator => "0011111101000000", --- 0.98828125 + j-0.152770996094
            im_multiplicator => "1111011000111001",
            data_re_out => mul_re_out(153),
            data_im_out => mul_im_out(153)
        );

 
    UMUL_154 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(154),
            data_im_in => first_stage_im_out(154),
            re_multiplicator => "0011111100110000", --- 0.9873046875 + j-0.158874511719
            im_multiplicator => "1111010111010101",
            data_re_out => mul_re_out(154),
            data_im_out => mul_im_out(154)
        );

 
    UMUL_155 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(155),
            data_im_in => first_stage_im_out(155),
            re_multiplicator => "0011111100100000", --- 0.986328125 + j-0.164916992188
            im_multiplicator => "1111010101110010",
            data_re_out => mul_re_out(155),
            data_im_out => mul_im_out(155)
        );

 
    UMUL_156 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(156),
            data_im_in => first_stage_im_out(156),
            re_multiplicator => "0011111100001111", --- 0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(156),
            data_im_out => mul_im_out(156)
        );

 
    UMUL_157 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(157),
            data_im_in => first_stage_im_out(157),
            re_multiplicator => "0011111011111101", --- 0.984191894531 + j-0.177001953125
            im_multiplicator => "1111010010101100",
            data_re_out => mul_re_out(157),
            data_im_out => mul_im_out(157)
        );

 
    UMUL_158 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(158),
            data_im_in => first_stage_im_out(158),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(158),
            data_im_out => mul_im_out(158)
        );

 
    UMUL_159 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(159),
            data_im_in => first_stage_im_out(159),
            re_multiplicator => "0011111011011000", --- 0.98193359375 + j-0.189086914062
            im_multiplicator => "1111001111100110",
            data_re_out => mul_re_out(159),
            data_im_out => mul_im_out(159)
        );

 
    UMUL_160 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(160),
            data_im_in => first_stage_im_out(160),
            re_multiplicator => "0011111011000101", --- 0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(160),
            data_im_out => mul_im_out(160)
        );

 
    UMUL_161 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(161),
            data_im_in => first_stage_im_out(161),
            re_multiplicator => "0011111010110001", --- 0.979553222656 + j-0.201110839844
            im_multiplicator => "1111001100100001",
            data_re_out => mul_re_out(161),
            data_im_out => mul_im_out(161)
        );

 
    UMUL_162 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(162),
            data_im_in => first_stage_im_out(162),
            re_multiplicator => "0011111010011101", --- 0.978332519531 + j-0.207092285156
            im_multiplicator => "1111001010111111",
            data_re_out => mul_re_out(162),
            data_im_out => mul_im_out(162)
        );

 
    UMUL_163 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(163),
            data_im_in => first_stage_im_out(163),
            re_multiplicator => "0011111010001000", --- 0.97705078125 + j-0.213134765625
            im_multiplicator => "1111001001011100",
            data_re_out => mul_re_out(163),
            data_im_out => mul_im_out(163)
        );

 
    UMUL_164 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(164),
            data_im_in => first_stage_im_out(164),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(164),
            data_im_out => mul_im_out(164)
        );

 
    UMUL_165 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(165),
            data_im_in => first_stage_im_out(165),
            re_multiplicator => "0011111001011100", --- 0.974365234375 + j-0.22509765625
            im_multiplicator => "1111000110011000",
            data_re_out => mul_re_out(165),
            data_im_out => mul_im_out(165)
        );

 
    UMUL_166 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(166),
            data_im_in => first_stage_im_out(166),
            re_multiplicator => "0011111001000101", --- 0.972961425781 + j-0.231079101562
            im_multiplicator => "1111000100110110",
            data_re_out => mul_re_out(166),
            data_im_out => mul_im_out(166)
        );

 
    UMUL_167 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(167),
            data_im_in => first_stage_im_out(167),
            re_multiplicator => "0011111000101101", --- 0.971496582031 + j-0.236999511719
            im_multiplicator => "1111000011010101",
            data_re_out => mul_re_out(167),
            data_im_out => mul_im_out(167)
        );

 
    UMUL_168 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(168),
            data_im_in => first_stage_im_out(168),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(168),
            data_im_out => mul_im_out(168)
        );

 
    UMUL_169 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(169),
            data_im_in => first_stage_im_out(169),
            re_multiplicator => "0011110111111100", --- 0.968505859375 + j-0.248901367188
            im_multiplicator => "1111000000010010",
            data_re_out => mul_re_out(169),
            data_im_out => mul_im_out(169)
        );

 
    UMUL_170 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(170),
            data_im_in => first_stage_im_out(170),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(170),
            data_im_out => mul_im_out(170)
        );

 
    UMUL_171 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(171),
            data_im_in => first_stage_im_out(171),
            re_multiplicator => "0011110111001001", --- 0.965393066406 + j-0.260803222656
            im_multiplicator => "1110111101001111",
            data_re_out => mul_re_out(171),
            data_im_out => mul_im_out(171)
        );

 
    UMUL_172 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(172),
            data_im_in => first_stage_im_out(172),
            re_multiplicator => "0011110110101111", --- 0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(172),
            data_im_out => mul_im_out(172)
        );

 
    UMUL_173 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(173),
            data_im_in => first_stage_im_out(173),
            re_multiplicator => "0011110110010011", --- 0.962097167969 + j-0.272644042969
            im_multiplicator => "1110111010001101",
            data_re_out => mul_re_out(173),
            data_im_out => mul_im_out(173)
        );

 
    UMUL_174 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(174),
            data_im_in => first_stage_im_out(174),
            re_multiplicator => "0011110101111000", --- 0.96044921875 + j-0.278503417969
            im_multiplicator => "1110111000101101",
            data_re_out => mul_re_out(174),
            data_im_out => mul_im_out(174)
        );

 
    UMUL_175 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(175),
            data_im_in => first_stage_im_out(175),
            re_multiplicator => "0011110101011011", --- 0.958679199219 + j-0.284423828125
            im_multiplicator => "1110110111001100",
            data_re_out => mul_re_out(175),
            data_im_out => mul_im_out(175)
        );

 
    UMUL_176 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(176),
            data_im_in => first_stage_im_out(176),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(176),
            data_im_out => mul_im_out(176)
        );

 
    UMUL_177 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(177),
            data_im_in => first_stage_im_out(177),
            re_multiplicator => "0011110100100001", --- 0.955139160156 + j-0.296142578125
            im_multiplicator => "1110110100001100",
            data_re_out => mul_re_out(177),
            data_im_out => mul_im_out(177)
        );

 
    UMUL_178 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(178),
            data_im_in => first_stage_im_out(178),
            re_multiplicator => "0011110100000011", --- 0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(178),
            data_im_out => mul_im_out(178)
        );

 
    UMUL_179 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(179),
            data_im_in => first_stage_im_out(179),
            re_multiplicator => "0011110011100100", --- 0.951416015625 + j-0.307861328125
            im_multiplicator => "1110110001001100",
            data_re_out => mul_re_out(179),
            data_im_out => mul_im_out(179)
        );

 
    UMUL_180 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(180),
            data_im_in => first_stage_im_out(180),
            re_multiplicator => "0011110011000101", --- 0.949523925781 + j-0.313659667969
            im_multiplicator => "1110101111101101",
            data_re_out => mul_re_out(180),
            data_im_out => mul_im_out(180)
        );

 
    UMUL_181 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(181),
            data_im_in => first_stage_im_out(181),
            re_multiplicator => "0011110010100101", --- 0.947570800781 + j-0.319519042969
            im_multiplicator => "1110101110001101",
            data_re_out => mul_re_out(181),
            data_im_out => mul_im_out(181)
        );

 
    UMUL_182 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(182),
            data_im_in => first_stage_im_out(182),
            re_multiplicator => "0011110010000101", --- 0.945617675781 + j-0.325317382812
            im_multiplicator => "1110101100101110",
            data_re_out => mul_re_out(182),
            data_im_out => mul_im_out(182)
        );

 
    UMUL_183 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(183),
            data_im_in => first_stage_im_out(183),
            re_multiplicator => "0011110001100100", --- 0.943603515625 + j-0.331115722656
            im_multiplicator => "1110101011001111",
            data_re_out => mul_re_out(183),
            data_im_out => mul_im_out(183)
        );

 
    UMUL_184 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(184),
            data_im_in => first_stage_im_out(184),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(184),
            data_im_out => mul_im_out(184)
        );

 
    UMUL_185 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(185),
            data_im_in => first_stage_im_out(185),
            re_multiplicator => "0011110000100000", --- 0.939453125 + j-0.342651367188
            im_multiplicator => "1110101000010010",
            data_re_out => mul_re_out(185),
            data_im_out => mul_im_out(185)
        );

 
    UMUL_186 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(186),
            data_im_in => first_stage_im_out(186),
            re_multiplicator => "0011101111111101", --- 0.937316894531 + j-0.348388671875
            im_multiplicator => "1110100110110100",
            data_re_out => mul_re_out(186),
            data_im_out => mul_im_out(186)
        );

 
    UMUL_187 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(187),
            data_im_in => first_stage_im_out(187),
            re_multiplicator => "0011101111011010", --- 0.935180664062 + j-0.354187011719
            im_multiplicator => "1110100101010101",
            data_re_out => mul_re_out(187),
            data_im_out => mul_im_out(187)
        );

 
    UMUL_188 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(188),
            data_im_in => first_stage_im_out(188),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(188),
            data_im_out => mul_im_out(188)
        );

 
    UMUL_189 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(189),
            data_im_in => first_stage_im_out(189),
            re_multiplicator => "0011101110010010", --- 0.930786132812 + j-0.365600585938
            im_multiplicator => "1110100010011010",
            data_re_out => mul_re_out(189),
            data_im_out => mul_im_out(189)
        );

 
    UMUL_190 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(190),
            data_im_in => first_stage_im_out(190),
            re_multiplicator => "0011101101101101", --- 0.928527832031 + j-0.371337890625
            im_multiplicator => "1110100000111100",
            data_re_out => mul_re_out(190),
            data_im_out => mul_im_out(190)
        );

 
    UMUL_191 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(191),
            data_im_in => first_stage_im_out(191),
            re_multiplicator => "0011101101000111", --- 0.926208496094 + j-0.377014160156
            im_multiplicator => "1110011111011111",
            data_re_out => mul_re_out(191),
            data_im_out => mul_im_out(191)
        );

 
    UMUL_192 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(192),
            data_im_in => first_stage_im_out(192),
            data_re_out => mul_re_out(192),
            data_im_out => mul_im_out(192)
        );

 
    UMUL_193 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(193),
            data_im_in => first_stage_im_out(193),
            re_multiplicator => "0011111111111111", --- 0.999938964844 + j-0.00921630859375
            im_multiplicator => "1111111101101001",
            data_re_out => mul_re_out(193),
            data_im_out => mul_im_out(193)
        );

 
    UMUL_194 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(194),
            data_im_in => first_stage_im_out(194),
            re_multiplicator => "0011111111111101", --- 0.999816894531 + j-0.0184326171875
            im_multiplicator => "1111111011010010",
            data_re_out => mul_re_out(194),
            data_im_out => mul_im_out(194)
        );

 
    UMUL_195 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(195),
            data_im_in => first_stage_im_out(195),
            re_multiplicator => "0011111111111010", --- 0.999633789062 + j-0.027587890625
            im_multiplicator => "1111111000111100",
            data_re_out => mul_re_out(195),
            data_im_out => mul_im_out(195)
        );

 
    UMUL_196 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(196),
            data_im_in => first_stage_im_out(196),
            re_multiplicator => "0011111111110101", --- 0.999328613281 + j-0.0368041992188
            im_multiplicator => "1111110110100101",
            data_re_out => mul_re_out(196),
            data_im_out => mul_im_out(196)
        );

 
    UMUL_197 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(197),
            data_im_in => first_stage_im_out(197),
            re_multiplicator => "0011111111101111", --- 0.998962402344 + j-0.0460205078125
            im_multiplicator => "1111110100001110",
            data_re_out => mul_re_out(197),
            data_im_out => mul_im_out(197)
        );

 
    UMUL_198 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(198),
            data_im_in => first_stage_im_out(198),
            re_multiplicator => "0011111111100111", --- 0.998474121094 + j-0.05517578125
            im_multiplicator => "1111110001111000",
            data_re_out => mul_re_out(198),
            data_im_out => mul_im_out(198)
        );

 
    UMUL_199 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(199),
            data_im_in => first_stage_im_out(199),
            re_multiplicator => "0011111111011110", --- 0.997924804688 + j-0.0643920898438
            im_multiplicator => "1111101111100001",
            data_re_out => mul_re_out(199),
            data_im_out => mul_im_out(199)
        );

 
    UMUL_200 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(200),
            data_im_in => first_stage_im_out(200),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(200),
            data_im_out => mul_im_out(200)
        );

 
    UMUL_201 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(201),
            data_im_in => first_stage_im_out(201),
            re_multiplicator => "0011111111001000", --- 0.99658203125 + j-0.082763671875
            im_multiplicator => "1111101010110100",
            data_re_out => mul_re_out(201),
            data_im_out => mul_im_out(201)
        );

 
    UMUL_202 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(202),
            data_im_in => first_stage_im_out(202),
            re_multiplicator => "0011111110111011", --- 0.995788574219 + j-0.0919189453125
            im_multiplicator => "1111101000011110",
            data_re_out => mul_re_out(202),
            data_im_out => mul_im_out(202)
        );

 
    UMUL_203 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(203),
            data_im_in => first_stage_im_out(203),
            re_multiplicator => "0011111110101100", --- 0.994873046875 + j-0.10107421875
            im_multiplicator => "1111100110001000",
            data_re_out => mul_re_out(203),
            data_im_out => mul_im_out(203)
        );

 
    UMUL_204 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(204),
            data_im_in => first_stage_im_out(204),
            re_multiplicator => "0011111110011100", --- 0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(204),
            data_im_out => mul_im_out(204)
        );

 
    UMUL_205 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(205),
            data_im_in => first_stage_im_out(205),
            re_multiplicator => "0011111110001011", --- 0.992858886719 + j-0.119384765625
            im_multiplicator => "1111100001011100",
            data_re_out => mul_re_out(205),
            data_im_out => mul_im_out(205)
        );

 
    UMUL_206 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(206),
            data_im_in => first_stage_im_out(206),
            re_multiplicator => "0011111101111000", --- 0.99169921875 + j-0.128479003906
            im_multiplicator => "1111011111000111",
            data_re_out => mul_re_out(206),
            data_im_out => mul_im_out(206)
        );

 
    UMUL_207 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(207),
            data_im_in => first_stage_im_out(207),
            re_multiplicator => "0011111101100100", --- 0.990478515625 + j-0.137634277344
            im_multiplicator => "1111011100110001",
            data_re_out => mul_re_out(207),
            data_im_out => mul_im_out(207)
        );

 
    UMUL_208 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(208),
            data_im_in => first_stage_im_out(208),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(208),
            data_im_out => mul_im_out(208)
        );

 
    UMUL_209 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(209),
            data_im_in => first_stage_im_out(209),
            re_multiplicator => "0011111100111000", --- 0.98779296875 + j-0.155822753906
            im_multiplicator => "1111011000000111",
            data_re_out => mul_re_out(209),
            data_im_out => mul_im_out(209)
        );

 
    UMUL_210 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(210),
            data_im_in => first_stage_im_out(210),
            re_multiplicator => "0011111100100000", --- 0.986328125 + j-0.164916992188
            im_multiplicator => "1111010101110010",
            data_re_out => mul_re_out(210),
            data_im_out => mul_im_out(210)
        );

 
    UMUL_211 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(211),
            data_im_in => first_stage_im_out(211),
            re_multiplicator => "0011111100000110", --- 0.984741210938 + j-0.174011230469
            im_multiplicator => "1111010011011101",
            data_re_out => mul_re_out(211),
            data_im_out => mul_im_out(211)
        );

 
    UMUL_212 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(212),
            data_im_in => first_stage_im_out(212),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(212),
            data_im_out => mul_im_out(212)
        );

 
    UMUL_213 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(213),
            data_im_in => first_stage_im_out(213),
            re_multiplicator => "0011111011001111", --- 0.981384277344 + j-0.192077636719
            im_multiplicator => "1111001110110101",
            data_re_out => mul_re_out(213),
            data_im_out => mul_im_out(213)
        );

 
    UMUL_214 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(214),
            data_im_in => first_stage_im_out(214),
            re_multiplicator => "0011111010110001", --- 0.979553222656 + j-0.201110839844
            im_multiplicator => "1111001100100001",
            data_re_out => mul_re_out(214),
            data_im_out => mul_im_out(214)
        );

 
    UMUL_215 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(215),
            data_im_in => first_stage_im_out(215),
            re_multiplicator => "0011111010010010", --- 0.977661132812 + j-0.210083007812
            im_multiplicator => "1111001010001110",
            data_re_out => mul_re_out(215),
            data_im_out => mul_im_out(215)
        );

 
    UMUL_216 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(216),
            data_im_in => first_stage_im_out(216),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(216),
            data_im_out => mul_im_out(216)
        );

 
    UMUL_217 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(217),
            data_im_in => first_stage_im_out(217),
            re_multiplicator => "0011111001010000", --- 0.9736328125 + j-0.228088378906
            im_multiplicator => "1111000101100111",
            data_re_out => mul_re_out(217),
            data_im_out => mul_im_out(217)
        );

 
    UMUL_218 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(218),
            data_im_in => first_stage_im_out(218),
            re_multiplicator => "0011111000101101", --- 0.971496582031 + j-0.236999511719
            im_multiplicator => "1111000011010101",
            data_re_out => mul_re_out(218),
            data_im_out => mul_im_out(218)
        );

 
    UMUL_219 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(219),
            data_im_in => first_stage_im_out(219),
            re_multiplicator => "0011111000001001", --- 0.969299316406 + j-0.245971679688
            im_multiplicator => "1111000001000010",
            data_re_out => mul_re_out(219),
            data_im_out => mul_im_out(219)
        );

 
    UMUL_220 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(220),
            data_im_in => first_stage_im_out(220),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(220),
            data_im_out => mul_im_out(220)
        );

 
    UMUL_221 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(221),
            data_im_in => first_stage_im_out(221),
            re_multiplicator => "0011110110111100", --- 0.964599609375 + j-0.263732910156
            im_multiplicator => "1110111100011111",
            data_re_out => mul_re_out(221),
            data_im_out => mul_im_out(221)
        );

 
    UMUL_222 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(222),
            data_im_in => first_stage_im_out(222),
            re_multiplicator => "0011110110010011", --- 0.962097167969 + j-0.272644042969
            im_multiplicator => "1110111010001101",
            data_re_out => mul_re_out(222),
            data_im_out => mul_im_out(222)
        );

 
    UMUL_223 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(223),
            data_im_in => first_stage_im_out(223),
            re_multiplicator => "0011110101101010", --- 0.959594726562 + j-0.281494140625
            im_multiplicator => "1110110111111100",
            data_re_out => mul_re_out(223),
            data_im_out => mul_im_out(223)
        );

 
    UMUL_224 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(224),
            data_im_in => first_stage_im_out(224),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(224),
            data_im_out => mul_im_out(224)
        );

 
    UMUL_225 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(225),
            data_im_in => first_stage_im_out(225),
            re_multiplicator => "0011110100010010", --- 0.954223632812 + j-0.299072265625
            im_multiplicator => "1110110011011100",
            data_re_out => mul_re_out(225),
            data_im_out => mul_im_out(225)
        );

 
    UMUL_226 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(226),
            data_im_in => first_stage_im_out(226),
            re_multiplicator => "0011110011100100", --- 0.951416015625 + j-0.307861328125
            im_multiplicator => "1110110001001100",
            data_re_out => mul_re_out(226),
            data_im_out => mul_im_out(226)
        );

 
    UMUL_227 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(227),
            data_im_in => first_stage_im_out(227),
            re_multiplicator => "0011110010110101", --- 0.948547363281 + j-0.316589355469
            im_multiplicator => "1110101110111101",
            data_re_out => mul_re_out(227),
            data_im_out => mul_im_out(227)
        );

 
    UMUL_228 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(228),
            data_im_in => first_stage_im_out(228),
            re_multiplicator => "0011110010000101", --- 0.945617675781 + j-0.325317382812
            im_multiplicator => "1110101100101110",
            data_re_out => mul_re_out(228),
            data_im_out => mul_im_out(228)
        );

 
    UMUL_229 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(229),
            data_im_in => first_stage_im_out(229),
            re_multiplicator => "0011110001010011", --- 0.942565917969 + j-0.333984375
            im_multiplicator => "1110101010100000",
            data_re_out => mul_re_out(229),
            data_im_out => mul_im_out(229)
        );

 
    UMUL_230 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(230),
            data_im_in => first_stage_im_out(230),
            re_multiplicator => "0011110000100000", --- 0.939453125 + j-0.342651367188
            im_multiplicator => "1110101000010010",
            data_re_out => mul_re_out(230),
            data_im_out => mul_im_out(230)
        );

 
    UMUL_231 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(231),
            data_im_in => first_stage_im_out(231),
            re_multiplicator => "0011101111101100", --- 0.936279296875 + j-0.351318359375
            im_multiplicator => "1110100110000100",
            data_re_out => mul_re_out(231),
            data_im_out => mul_im_out(231)
        );

 
    UMUL_232 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(232),
            data_im_in => first_stage_im_out(232),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(232),
            data_im_out => mul_im_out(232)
        );

 
    UMUL_233 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(233),
            data_im_in => first_stage_im_out(233),
            re_multiplicator => "0011101101111111", --- 0.929626464844 + j-0.368469238281
            im_multiplicator => "1110100001101011",
            data_re_out => mul_re_out(233),
            data_im_out => mul_im_out(233)
        );

 
    UMUL_234 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(234),
            data_im_in => first_stage_im_out(234),
            re_multiplicator => "0011101101000111", --- 0.926208496094 + j-0.377014160156
            im_multiplicator => "1110011111011111",
            data_re_out => mul_re_out(234),
            data_im_out => mul_im_out(234)
        );

 
    UMUL_235 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(235),
            data_im_in => first_stage_im_out(235),
            re_multiplicator => "0011101100001110", --- 0.922729492188 + j-0.385498046875
            im_multiplicator => "1110011101010100",
            data_re_out => mul_re_out(235),
            data_im_out => mul_im_out(235)
        );

 
    UMUL_236 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(236),
            data_im_in => first_stage_im_out(236),
            re_multiplicator => "0011101011010011", --- 0.919128417969 + j-0.393981933594
            im_multiplicator => "1110011011001001",
            data_re_out => mul_re_out(236),
            data_im_out => mul_im_out(236)
        );

 
    UMUL_237 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(237),
            data_im_in => first_stage_im_out(237),
            re_multiplicator => "0011101010010111", --- 0.915466308594 + j-0.402404785156
            im_multiplicator => "1110011000111111",
            data_re_out => mul_re_out(237),
            data_im_out => mul_im_out(237)
        );

 
    UMUL_238 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(238),
            data_im_in => first_stage_im_out(238),
            re_multiplicator => "0011101001011001", --- 0.911682128906 + j-0.410827636719
            im_multiplicator => "1110010110110101",
            data_re_out => mul_re_out(238),
            data_im_out => mul_im_out(238)
        );

 
    UMUL_239 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(239),
            data_im_in => first_stage_im_out(239),
            re_multiplicator => "0011101000011011", --- 0.907897949219 + j-0.419189453125
            im_multiplicator => "1110010100101100",
            data_re_out => mul_re_out(239),
            data_im_out => mul_im_out(239)
        );

 
    UMUL_240 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(240),
            data_im_in => first_stage_im_out(240),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(240),
            data_im_out => mul_im_out(240)
        );

 
    UMUL_241 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(241),
            data_im_in => first_stage_im_out(241),
            re_multiplicator => "0011100110011010", --- 0.900024414062 + j-0.435852050781
            im_multiplicator => "1110010000011011",
            data_re_out => mul_re_out(241),
            data_im_out => mul_im_out(241)
        );

 
    UMUL_242 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(242),
            data_im_in => first_stage_im_out(242),
            re_multiplicator => "0011100101011000", --- 0.89599609375 + j-0.444091796875
            im_multiplicator => "1110001110010100",
            data_re_out => mul_re_out(242),
            data_im_out => mul_im_out(242)
        );

 
    UMUL_243 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(243),
            data_im_in => first_stage_im_out(243),
            re_multiplicator => "0011100100010100", --- 0.891845703125 + j-0.452331542969
            im_multiplicator => "1110001100001101",
            data_re_out => mul_re_out(243),
            data_im_out => mul_im_out(243)
        );

 
    UMUL_244 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(244),
            data_im_in => first_stage_im_out(244),
            re_multiplicator => "0011100011001111", --- 0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(244),
            data_im_out => mul_im_out(244)
        );

 
    UMUL_245 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(245),
            data_im_in => first_stage_im_out(245),
            re_multiplicator => "0011100010001001", --- 0.883361816406 + j-0.468688964844
            im_multiplicator => "1110001000000001",
            data_re_out => mul_re_out(245),
            data_im_out => mul_im_out(245)
        );

 
    UMUL_246 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(246),
            data_im_in => first_stage_im_out(246),
            re_multiplicator => "0011100001000010", --- 0.879028320312 + j-0.476806640625
            im_multiplicator => "1110000101111100",
            data_re_out => mul_re_out(246),
            data_im_out => mul_im_out(246)
        );

 
    UMUL_247 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(247),
            data_im_in => first_stage_im_out(247),
            re_multiplicator => "0011011111111001", --- 0.874572753906 + j-0.48486328125
            im_multiplicator => "1110000011111000",
            data_re_out => mul_re_out(247),
            data_im_out => mul_im_out(247)
        );

 
    UMUL_248 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(248),
            data_im_in => first_stage_im_out(248),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(248),
            data_im_out => mul_im_out(248)
        );

 
    UMUL_249 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(249),
            data_im_in => first_stage_im_out(249),
            re_multiplicator => "0011011101100101", --- 0.865539550781 + j-0.500915527344
            im_multiplicator => "1101111111110001",
            data_re_out => mul_re_out(249),
            data_im_out => mul_im_out(249)
        );

 
    UMUL_250 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(250),
            data_im_in => first_stage_im_out(250),
            re_multiplicator => "0011011100011000", --- 0.86083984375 + j-0.508850097656
            im_multiplicator => "1101111101101111",
            data_re_out => mul_re_out(250),
            data_im_out => mul_im_out(250)
        );

 
    UMUL_251 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(251),
            data_im_in => first_stage_im_out(251),
            re_multiplicator => "0011011011001011", --- 0.856140136719 + j-0.516723632812
            im_multiplicator => "1101111011101110",
            data_re_out => mul_re_out(251),
            data_im_out => mul_im_out(251)
        );

 
    UMUL_252 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(252),
            data_im_in => first_stage_im_out(252),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(252),
            data_im_out => mul_im_out(252)
        );

 
    UMUL_253 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(253),
            data_im_in => first_stage_im_out(253),
            re_multiplicator => "0011011000101101", --- 0.846496582031 + j-0.532409667969
            im_multiplicator => "1101110111101101",
            data_re_out => mul_re_out(253),
            data_im_out => mul_im_out(253)
        );

 
    UMUL_254 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(254),
            data_im_in => first_stage_im_out(254),
            re_multiplicator => "0011010111011100", --- 0.841552734375 + j-0.540161132812
            im_multiplicator => "1101110101101110",
            data_re_out => mul_re_out(254),
            data_im_out => mul_im_out(254)
        );

 
    UMUL_255 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(255),
            data_im_in => first_stage_im_out(255),
            re_multiplicator => "0011010110001010", --- 0.836547851562 + j-0.547912597656
            im_multiplicator => "1101110011101111",
            data_re_out => mul_re_out(255),
            data_im_out => mul_im_out(255)
        );

 
    UMUL_256 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(256),
            data_im_in => first_stage_im_out(256),
            data_re_out => mul_re_out(256),
            data_im_out => mul_im_out(256)
        );

 
    UMUL_257 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(257),
            data_im_in => first_stage_im_out(257),
            re_multiplicator => "0011111111111111", --- 0.999938964844 + j-0.0122680664062
            im_multiplicator => "1111111100110111",
            data_re_out => mul_re_out(257),
            data_im_out => mul_im_out(257)
        );

 
    UMUL_258 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(258),
            data_im_in => first_stage_im_out(258),
            re_multiplicator => "0011111111111011", --- 0.999694824219 + j-0.0245361328125
            im_multiplicator => "1111111001101110",
            data_re_out => mul_re_out(258),
            data_im_out => mul_im_out(258)
        );

 
    UMUL_259 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(259),
            data_im_in => first_stage_im_out(259),
            re_multiplicator => "0011111111110101", --- 0.999328613281 + j-0.0368041992188
            im_multiplicator => "1111110110100101",
            data_re_out => mul_re_out(259),
            data_im_out => mul_im_out(259)
        );

 
    UMUL_260 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(260),
            data_im_in => first_stage_im_out(260),
            re_multiplicator => "0011111111101100", --- 0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(260),
            data_im_out => mul_im_out(260)
        );

 
    UMUL_261 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(261),
            data_im_in => first_stage_im_out(261),
            re_multiplicator => "0011111111100001", --- 0.998107910156 + j-0.0613403320312
            im_multiplicator => "1111110000010011",
            data_re_out => mul_re_out(261),
            data_im_out => mul_im_out(261)
        );

 
    UMUL_262 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(262),
            data_im_in => first_stage_im_out(262),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(262),
            data_im_out => mul_im_out(262)
        );

 
    UMUL_263 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(263),
            data_im_in => first_stage_im_out(263),
            re_multiplicator => "0011111111000100", --- 0.996337890625 + j-0.0858154296875
            im_multiplicator => "1111101010000010",
            data_re_out => mul_re_out(263),
            data_im_out => mul_im_out(263)
        );

 
    UMUL_264 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(264),
            data_im_in => first_stage_im_out(264),
            re_multiplicator => "0011111110110001", --- 0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(264),
            data_im_out => mul_im_out(264)
        );

 
    UMUL_265 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(265),
            data_im_in => first_stage_im_out(265),
            re_multiplicator => "0011111110011100", --- 0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(265),
            data_im_out => mul_im_out(265)
        );

 
    UMUL_266 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(266),
            data_im_in => first_stage_im_out(266),
            re_multiplicator => "0011111110000101", --- 0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(266),
            data_im_out => mul_im_out(266)
        );

 
    UMUL_267 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(267),
            data_im_in => first_stage_im_out(267),
            re_multiplicator => "0011111101101011", --- 0.990905761719 + j-0.134582519531
            im_multiplicator => "1111011101100011",
            data_re_out => mul_re_out(267),
            data_im_out => mul_im_out(267)
        );

 
    UMUL_268 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(268),
            data_im_in => first_stage_im_out(268),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(268),
            data_im_out => mul_im_out(268)
        );

 
    UMUL_269 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(269),
            data_im_in => first_stage_im_out(269),
            re_multiplicator => "0011111100110000", --- 0.9873046875 + j-0.158874511719
            im_multiplicator => "1111010111010101",
            data_re_out => mul_re_out(269),
            data_im_out => mul_im_out(269)
        );

 
    UMUL_270 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(270),
            data_im_in => first_stage_im_out(270),
            re_multiplicator => "0011111100001111", --- 0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(270),
            data_im_out => mul_im_out(270)
        );

 
    UMUL_271 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(271),
            data_im_in => first_stage_im_out(271),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(271),
            data_im_out => mul_im_out(271)
        );

 
    UMUL_272 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(272),
            data_im_in => first_stage_im_out(272),
            re_multiplicator => "0011111011000101", --- 0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(272),
            data_im_out => mul_im_out(272)
        );

 
    UMUL_273 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(273),
            data_im_in => first_stage_im_out(273),
            re_multiplicator => "0011111010011101", --- 0.978332519531 + j-0.207092285156
            im_multiplicator => "1111001010111111",
            data_re_out => mul_re_out(273),
            data_im_out => mul_im_out(273)
        );

 
    UMUL_274 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(274),
            data_im_in => first_stage_im_out(274),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(274),
            data_im_out => mul_im_out(274)
        );

 
    UMUL_275 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(275),
            data_im_in => first_stage_im_out(275),
            re_multiplicator => "0011111001000101", --- 0.972961425781 + j-0.231079101562
            im_multiplicator => "1111000100110110",
            data_re_out => mul_re_out(275),
            data_im_out => mul_im_out(275)
        );

 
    UMUL_276 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(276),
            data_im_in => first_stage_im_out(276),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(276),
            data_im_out => mul_im_out(276)
        );

 
    UMUL_277 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(277),
            data_im_in => first_stage_im_out(277),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(277),
            data_im_out => mul_im_out(277)
        );

 
    UMUL_278 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(278),
            data_im_in => first_stage_im_out(278),
            re_multiplicator => "0011110110101111", --- 0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(278),
            data_im_out => mul_im_out(278)
        );

 
    UMUL_279 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(279),
            data_im_in => first_stage_im_out(279),
            re_multiplicator => "0011110101111000", --- 0.96044921875 + j-0.278503417969
            im_multiplicator => "1110111000101101",
            data_re_out => mul_re_out(279),
            data_im_out => mul_im_out(279)
        );

 
    UMUL_280 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(280),
            data_im_in => first_stage_im_out(280),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(280),
            data_im_out => mul_im_out(280)
        );

 
    UMUL_281 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(281),
            data_im_in => first_stage_im_out(281),
            re_multiplicator => "0011110100000011", --- 0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(281),
            data_im_out => mul_im_out(281)
        );

 
    UMUL_282 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(282),
            data_im_in => first_stage_im_out(282),
            re_multiplicator => "0011110011000101", --- 0.949523925781 + j-0.313659667969
            im_multiplicator => "1110101111101101",
            data_re_out => mul_re_out(282),
            data_im_out => mul_im_out(282)
        );

 
    UMUL_283 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(283),
            data_im_in => first_stage_im_out(283),
            re_multiplicator => "0011110010000101", --- 0.945617675781 + j-0.325317382812
            im_multiplicator => "1110101100101110",
            data_re_out => mul_re_out(283),
            data_im_out => mul_im_out(283)
        );

 
    UMUL_284 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(284),
            data_im_in => first_stage_im_out(284),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(284),
            data_im_out => mul_im_out(284)
        );

 
    UMUL_285 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(285),
            data_im_in => first_stage_im_out(285),
            re_multiplicator => "0011101111111101", --- 0.937316894531 + j-0.348388671875
            im_multiplicator => "1110100110110100",
            data_re_out => mul_re_out(285),
            data_im_out => mul_im_out(285)
        );

 
    UMUL_286 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(286),
            data_im_in => first_stage_im_out(286),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(286),
            data_im_out => mul_im_out(286)
        );

 
    UMUL_287 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(287),
            data_im_in => first_stage_im_out(287),
            re_multiplicator => "0011101101101101", --- 0.928527832031 + j-0.371337890625
            im_multiplicator => "1110100000111100",
            data_re_out => mul_re_out(287),
            data_im_out => mul_im_out(287)
        );

 
    UMUL_288 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(288),
            data_im_in => first_stage_im_out(288),
            re_multiplicator => "0011101100100001", --- 0.923889160156 + j-0.382690429688
            im_multiplicator => "1110011110000010",
            data_re_out => mul_re_out(288),
            data_im_out => mul_im_out(288)
        );

 
    UMUL_289 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(289),
            data_im_in => first_stage_im_out(289),
            re_multiplicator => "0011101011010011", --- 0.919128417969 + j-0.393981933594
            im_multiplicator => "1110011011001001",
            data_re_out => mul_re_out(289),
            data_im_out => mul_im_out(289)
        );

 
    UMUL_290 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(290),
            data_im_in => first_stage_im_out(290),
            re_multiplicator => "0011101010000010", --- 0.914184570312 + j-0.405212402344
            im_multiplicator => "1110011000010001",
            data_re_out => mul_re_out(290),
            data_im_out => mul_im_out(290)
        );

 
    UMUL_291 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(291),
            data_im_in => first_stage_im_out(291),
            re_multiplicator => "0011101000110000", --- 0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(291),
            data_im_out => mul_im_out(291)
        );

 
    UMUL_292 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(292),
            data_im_in => first_stage_im_out(292),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(292),
            data_im_out => mul_im_out(292)
        );

 
    UMUL_293 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(293),
            data_im_in => first_stage_im_out(293),
            re_multiplicator => "0011100110000100", --- 0.898681640625 + j-0.438598632812
            im_multiplicator => "1110001111101110",
            data_re_out => mul_re_out(293),
            data_im_out => mul_im_out(293)
        );

 
    UMUL_294 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(294),
            data_im_in => first_stage_im_out(294),
            re_multiplicator => "0011100100101011", --- 0.893249511719 + j-0.449584960938
            im_multiplicator => "1110001100111010",
            data_re_out => mul_re_out(294),
            data_im_out => mul_im_out(294)
        );

 
    UMUL_295 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(295),
            data_im_in => first_stage_im_out(295),
            re_multiplicator => "0011100011001111", --- 0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(295),
            data_im_out => mul_im_out(295)
        );

 
    UMUL_296 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(296),
            data_im_in => first_stage_im_out(296),
            re_multiplicator => "0011100001110001", --- 0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(296),
            data_im_out => mul_im_out(296)
        );

 
    UMUL_297 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(297),
            data_im_in => first_stage_im_out(297),
            re_multiplicator => "0011100000010010", --- 0.876098632812 + j-0.482177734375
            im_multiplicator => "1110000100100100",
            data_re_out => mul_re_out(297),
            data_im_out => mul_im_out(297)
        );

 
    UMUL_298 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(298),
            data_im_in => first_stage_im_out(298),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(298),
            data_im_out => mul_im_out(298)
        );

 
    UMUL_299 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(299),
            data_im_in => first_stage_im_out(299),
            re_multiplicator => "0011011101001011", --- 0.863952636719 + j-0.503540039062
            im_multiplicator => "1101111111000110",
            data_re_out => mul_re_out(299),
            data_im_out => mul_im_out(299)
        );

 
    UMUL_300 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(300),
            data_im_in => first_stage_im_out(300),
            re_multiplicator => "0011011011100101", --- 0.857727050781 + j-0.514099121094
            im_multiplicator => "1101111100011001",
            data_re_out => mul_re_out(300),
            data_im_out => mul_im_out(300)
        );

 
    UMUL_301 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(301),
            data_im_in => first_stage_im_out(301),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(301),
            data_im_out => mul_im_out(301)
        );

 
    UMUL_302 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(302),
            data_im_in => first_stage_im_out(302),
            re_multiplicator => "0011011000010010", --- 0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(302),
            data_im_out => mul_im_out(302)
        );

 
    UMUL_303 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(303),
            data_im_in => first_stage_im_out(303),
            re_multiplicator => "0011010110100101", --- 0.838195800781 + j-0.545349121094
            im_multiplicator => "1101110100011001",
            data_re_out => mul_re_out(303),
            data_im_out => mul_im_out(303)
        );

 
    UMUL_304 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(304),
            data_im_in => first_stage_im_out(304),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(304),
            data_im_out => mul_im_out(304)
        );

 
    UMUL_305 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(305),
            data_im_in => first_stage_im_out(305),
            re_multiplicator => "0011010011000110", --- 0.824584960938 + j-0.565734863281
            im_multiplicator => "1101101111001011",
            data_re_out => mul_re_out(305),
            data_im_out => mul_im_out(305)
        );

 
    UMUL_306 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(306),
            data_im_in => first_stage_im_out(306),
            re_multiplicator => "0011010001010011", --- 0.817565917969 + j-0.575805664062
            im_multiplicator => "1101101100100110",
            data_re_out => mul_re_out(306),
            data_im_out => mul_im_out(306)
        );

 
    UMUL_307 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(307),
            data_im_in => first_stage_im_out(307),
            re_multiplicator => "0011001111011111", --- 0.810485839844 + j-0.585815429688
            im_multiplicator => "1101101010000010",
            data_re_out => mul_re_out(307),
            data_im_out => mul_im_out(307)
        );

 
    UMUL_308 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(308),
            data_im_in => first_stage_im_out(308),
            re_multiplicator => "0011001101101000", --- 0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(308),
            data_im_out => mul_im_out(308)
        );

 
    UMUL_309 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(309),
            data_im_in => first_stage_im_out(309),
            re_multiplicator => "0011001011101111", --- 0.795837402344 + j-0.605529785156
            im_multiplicator => "1101100100111111",
            data_re_out => mul_re_out(309),
            data_im_out => mul_im_out(309)
        );

 
    UMUL_310 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(310),
            data_im_in => first_stage_im_out(310),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(310),
            data_im_out => mul_im_out(310)
        );

 
    UMUL_311 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(311),
            data_im_in => first_stage_im_out(311),
            re_multiplicator => "0011000111111000", --- 0.78076171875 + j-0.624877929688
            im_multiplicator => "1101100000000010",
            data_re_out => mul_re_out(311),
            data_im_out => mul_im_out(311)
        );

 
    UMUL_312 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(312),
            data_im_in => first_stage_im_out(312),
            re_multiplicator => "0011000101111001", --- 0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(312),
            data_im_out => mul_im_out(312)
        );

 
    UMUL_313 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(313),
            data_im_in => first_stage_im_out(313),
            re_multiplicator => "0011000011111001", --- 0.765197753906 + j-0.643859863281
            im_multiplicator => "1101011011001011",
            data_re_out => mul_re_out(313),
            data_im_out => mul_im_out(313)
        );

 
    UMUL_314 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(314),
            data_im_in => first_stage_im_out(314),
            re_multiplicator => "0011000001110110", --- 0.757202148438 + j-0.653198242188
            im_multiplicator => "1101011000110010",
            data_re_out => mul_re_out(314),
            data_im_out => mul_im_out(314)
        );

 
    UMUL_315 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(315),
            data_im_in => first_stage_im_out(315),
            re_multiplicator => "0010111111110010", --- 0.749145507812 + j-0.662414550781
            im_multiplicator => "1101010110011011",
            data_re_out => mul_re_out(315),
            data_im_out => mul_im_out(315)
        );

 
    UMUL_316 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(316),
            data_im_in => first_stage_im_out(316),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(316),
            data_im_out => mul_im_out(316)
        );

 
    UMUL_317 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(317),
            data_im_in => first_stage_im_out(317),
            re_multiplicator => "0010111011100100", --- 0.732666015625 + j-0.680603027344
            im_multiplicator => "1101010001110001",
            data_re_out => mul_re_out(317),
            data_im_out => mul_im_out(317)
        );

 
    UMUL_318 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(318),
            data_im_in => first_stage_im_out(318),
            re_multiplicator => "0010111001011010", --- 0.724243164062 + j-0.689514160156
            im_multiplicator => "1101001111011111",
            data_re_out => mul_re_out(318),
            data_im_out => mul_im_out(318)
        );

 
    UMUL_319 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(319),
            data_im_in => first_stage_im_out(319),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(319),
            data_im_out => mul_im_out(319)
        );

 
    UMUL_320 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(320),
            data_im_in => first_stage_im_out(320),
            data_re_out => mul_re_out(320),
            data_im_out => mul_im_out(320)
        );

 
    UMUL_321 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(321),
            data_im_in => first_stage_im_out(321),
            re_multiplicator => "0011111111111110", --- 0.999877929688 + j-0.0153198242188
            im_multiplicator => "1111111100000101",
            data_re_out => mul_re_out(321),
            data_im_out => mul_im_out(321)
        );

 
    UMUL_322 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(322),
            data_im_in => first_stage_im_out(322),
            re_multiplicator => "0011111111111000", --- 0.99951171875 + j-0.0307006835938
            im_multiplicator => "1111111000001001",
            data_re_out => mul_re_out(322),
            data_im_out => mul_im_out(322)
        );

 
    UMUL_323 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(323),
            data_im_in => first_stage_im_out(323),
            re_multiplicator => "0011111111101111", --- 0.998962402344 + j-0.0460205078125
            im_multiplicator => "1111110100001110",
            data_re_out => mul_re_out(323),
            data_im_out => mul_im_out(323)
        );

 
    UMUL_324 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(324),
            data_im_in => first_stage_im_out(324),
            re_multiplicator => "0011111111100001", --- 0.998107910156 + j-0.0613403320312
            im_multiplicator => "1111110000010011",
            data_re_out => mul_re_out(324),
            data_im_out => mul_im_out(324)
        );

 
    UMUL_325 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(325),
            data_im_in => first_stage_im_out(325),
            re_multiplicator => "0011111111010000", --- 0.9970703125 + j-0.0765991210938
            im_multiplicator => "1111101100011001",
            data_re_out => mul_re_out(325),
            data_im_out => mul_im_out(325)
        );

 
    UMUL_326 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(326),
            data_im_in => first_stage_im_out(326),
            re_multiplicator => "0011111110111011", --- 0.995788574219 + j-0.0919189453125
            im_multiplicator => "1111101000011110",
            data_re_out => mul_re_out(326),
            data_im_out => mul_im_out(326)
        );

 
    UMUL_327 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(327),
            data_im_in => first_stage_im_out(327),
            re_multiplicator => "0011111110100010", --- 0.994262695312 + j-0.107177734375
            im_multiplicator => "1111100100100100",
            data_re_out => mul_re_out(327),
            data_im_out => mul_im_out(327)
        );

 
    UMUL_328 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(328),
            data_im_in => first_stage_im_out(328),
            re_multiplicator => "0011111110000101", --- 0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(328),
            data_im_out => mul_im_out(328)
        );

 
    UMUL_329 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(329),
            data_im_in => first_stage_im_out(329),
            re_multiplicator => "0011111101100100", --- 0.990478515625 + j-0.137634277344
            im_multiplicator => "1111011100110001",
            data_re_out => mul_re_out(329),
            data_im_out => mul_im_out(329)
        );

 
    UMUL_330 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(330),
            data_im_in => first_stage_im_out(330),
            re_multiplicator => "0011111101000000", --- 0.98828125 + j-0.152770996094
            im_multiplicator => "1111011000111001",
            data_re_out => mul_re_out(330),
            data_im_out => mul_im_out(330)
        );

 
    UMUL_331 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(331),
            data_im_in => first_stage_im_out(331),
            re_multiplicator => "0011111100010111", --- 0.985778808594 + j-0.16796875
            im_multiplicator => "1111010101000000",
            data_re_out => mul_re_out(331),
            data_im_out => mul_im_out(331)
        );

 
    UMUL_332 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(332),
            data_im_in => first_stage_im_out(332),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(332),
            data_im_out => mul_im_out(332)
        );

 
    UMUL_333 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(333),
            data_im_in => first_stage_im_out(333),
            re_multiplicator => "0011111010111011", --- 0.980163574219 + j-0.198120117188
            im_multiplicator => "1111001101010010",
            data_re_out => mul_re_out(333),
            data_im_out => mul_im_out(333)
        );

 
    UMUL_334 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(334),
            data_im_in => first_stage_im_out(334),
            re_multiplicator => "0011111010001000", --- 0.97705078125 + j-0.213134765625
            im_multiplicator => "1111001001011100",
            data_re_out => mul_re_out(334),
            data_im_out => mul_im_out(334)
        );

 
    UMUL_335 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(335),
            data_im_in => first_stage_im_out(335),
            re_multiplicator => "0011111001010000", --- 0.9736328125 + j-0.228088378906
            im_multiplicator => "1111000101100111",
            data_re_out => mul_re_out(335),
            data_im_out => mul_im_out(335)
        );

 
    UMUL_336 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(336),
            data_im_in => first_stage_im_out(336),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(336),
            data_im_out => mul_im_out(336)
        );

 
    UMUL_337 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(337),
            data_im_in => first_stage_im_out(337),
            re_multiplicator => "0011110111010110", --- 0.966186523438 + j-0.2578125
            im_multiplicator => "1110111110000000",
            data_re_out => mul_re_out(337),
            data_im_out => mul_im_out(337)
        );

 
    UMUL_338 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(338),
            data_im_in => first_stage_im_out(338),
            re_multiplicator => "0011110110010011", --- 0.962097167969 + j-0.272644042969
            im_multiplicator => "1110111010001101",
            data_re_out => mul_re_out(338),
            data_im_out => mul_im_out(338)
        );

 
    UMUL_339 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(339),
            data_im_in => first_stage_im_out(339),
            re_multiplicator => "0011110101001101", --- 0.957824707031 + j-0.287353515625
            im_multiplicator => "1110110110011100",
            data_re_out => mul_re_out(339),
            data_im_out => mul_im_out(339)
        );

 
    UMUL_340 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(340),
            data_im_in => first_stage_im_out(340),
            re_multiplicator => "0011110100000011", --- 0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(340),
            data_im_out => mul_im_out(340)
        );

 
    UMUL_341 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(341),
            data_im_in => first_stage_im_out(341),
            re_multiplicator => "0011110010110101", --- 0.948547363281 + j-0.316589355469
            im_multiplicator => "1110101110111101",
            data_re_out => mul_re_out(341),
            data_im_out => mul_im_out(341)
        );

 
    UMUL_342 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(342),
            data_im_in => first_stage_im_out(342),
            re_multiplicator => "0011110001100100", --- 0.943603515625 + j-0.331115722656
            im_multiplicator => "1110101011001111",
            data_re_out => mul_re_out(342),
            data_im_out => mul_im_out(342)
        );

 
    UMUL_343 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(343),
            data_im_in => first_stage_im_out(343),
            re_multiplicator => "0011110000001111", --- 0.938415527344 + j-0.345520019531
            im_multiplicator => "1110100111100011",
            data_re_out => mul_re_out(343),
            data_im_out => mul_im_out(343)
        );

 
    UMUL_344 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(344),
            data_im_in => first_stage_im_out(344),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(344),
            data_im_out => mul_im_out(344)
        );

 
    UMUL_345 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(345),
            data_im_in => first_stage_im_out(345),
            re_multiplicator => "0011101101011010", --- 0.927368164062 + j-0.374145507812
            im_multiplicator => "1110100000001110",
            data_re_out => mul_re_out(345),
            data_im_out => mul_im_out(345)
        );

 
    UMUL_346 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(346),
            data_im_in => first_stage_im_out(346),
            re_multiplicator => "0011101011111010", --- 0.921508789062 + j-0.388366699219
            im_multiplicator => "1110011100100101",
            data_re_out => mul_re_out(346),
            data_im_out => mul_im_out(346)
        );

 
    UMUL_347 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(347),
            data_im_in => first_stage_im_out(347),
            re_multiplicator => "0011101010010111", --- 0.915466308594 + j-0.402404785156
            im_multiplicator => "1110011000111111",
            data_re_out => mul_re_out(347),
            data_im_out => mul_im_out(347)
        );

 
    UMUL_348 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(348),
            data_im_in => first_stage_im_out(348),
            re_multiplicator => "0011101000110000", --- 0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(348),
            data_im_out => mul_im_out(348)
        );

 
    UMUL_349 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(349),
            data_im_in => first_stage_im_out(349),
            re_multiplicator => "0011100111000101", --- 0.902648925781 + j-0.430297851562
            im_multiplicator => "1110010001110110",
            data_re_out => mul_re_out(349),
            data_im_out => mul_im_out(349)
        );

 
    UMUL_350 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(350),
            data_im_in => first_stage_im_out(350),
            re_multiplicator => "0011100101011000", --- 0.89599609375 + j-0.444091796875
            im_multiplicator => "1110001110010100",
            data_re_out => mul_re_out(350),
            data_im_out => mul_im_out(350)
        );

 
    UMUL_351 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(351),
            data_im_in => first_stage_im_out(351),
            re_multiplicator => "0011100011100110", --- 0.889038085938 + j-0.457824707031
            im_multiplicator => "1110001010110011",
            data_re_out => mul_re_out(351),
            data_im_out => mul_im_out(351)
        );

 
    UMUL_352 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(352),
            data_im_in => first_stage_im_out(352),
            re_multiplicator => "0011100001110001", --- 0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(352),
            data_im_out => mul_im_out(352)
        );

 
    UMUL_353 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(353),
            data_im_in => first_stage_im_out(353),
            re_multiplicator => "0011011111111001", --- 0.874572753906 + j-0.48486328125
            im_multiplicator => "1110000011111000",
            data_re_out => mul_re_out(353),
            data_im_out => mul_im_out(353)
        );

 
    UMUL_354 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(354),
            data_im_in => first_stage_im_out(354),
            re_multiplicator => "0011011101111110", --- 0.867065429688 + j-0.498229980469
            im_multiplicator => "1110000000011101",
            data_re_out => mul_re_out(354),
            data_im_out => mul_im_out(354)
        );

 
    UMUL_355 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(355),
            data_im_in => first_stage_im_out(355),
            re_multiplicator => "0011011011111111", --- 0.859313964844 + j-0.511474609375
            im_multiplicator => "1101111101000100",
            data_re_out => mul_re_out(355),
            data_im_out => mul_im_out(355)
        );

 
    UMUL_356 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(356),
            data_im_in => first_stage_im_out(356),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(356),
            data_im_out => mul_im_out(356)
        );

 
    UMUL_357 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(357),
            data_im_in => first_stage_im_out(357),
            re_multiplicator => "0011010111110111", --- 0.843200683594 + j-0.53759765625
            im_multiplicator => "1101110110011000",
            data_re_out => mul_re_out(357),
            data_im_out => mul_im_out(357)
        );

 
    UMUL_358 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(358),
            data_im_in => first_stage_im_out(358),
            re_multiplicator => "0011010101101110", --- 0.834838867188 + j-0.550476074219
            im_multiplicator => "1101110011000101",
            data_re_out => mul_re_out(358),
            data_im_out => mul_im_out(358)
        );

 
    UMUL_359 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(359),
            data_im_in => first_stage_im_out(359),
            re_multiplicator => "0011010011100010", --- 0.826293945312 + j-0.563171386719
            im_multiplicator => "1101101111110101",
            data_re_out => mul_re_out(359),
            data_im_out => mul_im_out(359)
        );

 
    UMUL_360 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(360),
            data_im_in => first_stage_im_out(360),
            re_multiplicator => "0011010001010011", --- 0.817565917969 + j-0.575805664062
            im_multiplicator => "1101101100100110",
            data_re_out => mul_re_out(360),
            data_im_out => mul_im_out(360)
        );

 
    UMUL_361 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(361),
            data_im_in => first_stage_im_out(361),
            re_multiplicator => "0011001111000001", --- 0.808654785156 + j-0.588256835938
            im_multiplicator => "1101101001011010",
            data_re_out => mul_re_out(361),
            data_im_out => mul_im_out(361)
        );

 
    UMUL_362 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(362),
            data_im_in => first_stage_im_out(362),
            re_multiplicator => "0011001100101100", --- 0.799560546875 + j-0.600646972656
            im_multiplicator => "1101100110001111",
            data_re_out => mul_re_out(362),
            data_im_out => mul_im_out(362)
        );

 
    UMUL_363 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(363),
            data_im_in => first_stage_im_out(363),
            re_multiplicator => "0011001010010011", --- 0.790222167969 + j-0.61279296875
            im_multiplicator => "1101100011001000",
            data_re_out => mul_re_out(363),
            data_im_out => mul_im_out(363)
        );

 
    UMUL_364 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(364),
            data_im_in => first_stage_im_out(364),
            re_multiplicator => "0011000111111000", --- 0.78076171875 + j-0.624877929688
            im_multiplicator => "1101100000000010",
            data_re_out => mul_re_out(364),
            data_im_out => mul_im_out(364)
        );

 
    UMUL_365 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(365),
            data_im_in => first_stage_im_out(365),
            re_multiplicator => "0011000101011001", --- 0.771057128906 + j-0.636779785156
            im_multiplicator => "1101011100111111",
            data_re_out => mul_re_out(365),
            data_im_out => mul_im_out(365)
        );

 
    UMUL_366 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(366),
            data_im_in => first_stage_im_out(366),
            re_multiplicator => "0011000010111000", --- 0.76123046875 + j-0.648498535156
            im_multiplicator => "1101011001111111",
            data_re_out => mul_re_out(366),
            data_im_out => mul_im_out(366)
        );

 
    UMUL_367 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(367),
            data_im_in => first_stage_im_out(367),
            re_multiplicator => "0011000000010011", --- 0.751159667969 + j-0.660095214844
            im_multiplicator => "1101010111000001",
            data_re_out => mul_re_out(367),
            data_im_out => mul_im_out(367)
        );

 
    UMUL_368 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(368),
            data_im_in => first_stage_im_out(368),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(368),
            data_im_out => mul_im_out(368)
        );

 
    UMUL_369 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(369),
            data_im_in => first_stage_im_out(369),
            re_multiplicator => "0010111011000010", --- 0.730590820312 + j-0.682861328125
            im_multiplicator => "1101010001001100",
            data_re_out => mul_re_out(369),
            data_im_out => mul_im_out(369)
        );

 
    UMUL_370 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(370),
            data_im_in => first_stage_im_out(370),
            re_multiplicator => "0010111000010101", --- 0.720031738281 + j-0.693969726562
            im_multiplicator => "1101001110010110",
            data_re_out => mul_re_out(370),
            data_im_out => mul_im_out(370)
        );

 
    UMUL_371 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(371),
            data_im_in => first_stage_im_out(371),
            re_multiplicator => "0010110101100101", --- 0.709289550781 + j-0.704956054688
            im_multiplicator => "1101001011100010",
            data_re_out => mul_re_out(371),
            data_im_out => mul_im_out(371)
        );

 
    UMUL_372 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(372),
            data_im_in => first_stage_im_out(372),
            re_multiplicator => "0010110010110010", --- 0.698364257812 + j-0.715759277344
            im_multiplicator => "1101001000110001",
            data_re_out => mul_re_out(372),
            data_im_out => mul_im_out(372)
        );

 
    UMUL_373 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(373),
            data_im_in => first_stage_im_out(373),
            re_multiplicator => "0010101111111101", --- 0.687316894531 + j-0.726379394531
            im_multiplicator => "1101000110000011",
            data_re_out => mul_re_out(373),
            data_im_out => mul_im_out(373)
        );

 
    UMUL_374 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(374),
            data_im_in => first_stage_im_out(374),
            re_multiplicator => "0010101101000101", --- 0.676086425781 + j-0.73681640625
            im_multiplicator => "1101000011011000",
            data_re_out => mul_re_out(374),
            data_im_out => mul_im_out(374)
        );

 
    UMUL_375 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(375),
            data_im_in => first_stage_im_out(375),
            re_multiplicator => "0010101010001011", --- 0.664733886719 + j-0.7470703125
            im_multiplicator => "1101000000110000",
            data_re_out => mul_re_out(375),
            data_im_out => mul_im_out(375)
        );

 
    UMUL_376 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(376),
            data_im_in => first_stage_im_out(376),
            re_multiplicator => "0010100111001110", --- 0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(376),
            data_im_out => mul_im_out(376)
        );

 
    UMUL_377 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(377),
            data_im_in => first_stage_im_out(377),
            re_multiplicator => "0010100100001110", --- 0.641479492188 + j-0.767150878906
            im_multiplicator => "1100111011100111",
            data_re_out => mul_re_out(377),
            data_im_out => mul_im_out(377)
        );

 
    UMUL_378 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(378),
            data_im_in => first_stage_im_out(378),
            re_multiplicator => "0010100001001100", --- 0.629638671875 + j-0.776916503906
            im_multiplicator => "1100111001000111",
            data_re_out => mul_re_out(378),
            data_im_out => mul_im_out(378)
        );

 
    UMUL_379 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(379),
            data_im_in => first_stage_im_out(379),
            re_multiplicator => "0010011110001000", --- 0.61767578125 + j-0.786437988281
            im_multiplicator => "1100110110101011",
            data_re_out => mul_re_out(379),
            data_im_out => mul_im_out(379)
        );

 
    UMUL_380 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(380),
            data_im_in => first_stage_im_out(380),
            re_multiplicator => "0010011011000001", --- 0.605529785156 + j-0.795837402344
            im_multiplicator => "1100110100010001",
            data_re_out => mul_re_out(380),
            data_im_out => mul_im_out(380)
        );

 
    UMUL_381 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(381),
            data_im_in => first_stage_im_out(381),
            re_multiplicator => "0010010111111000", --- 0.59326171875 + j-0.805053710938
            im_multiplicator => "1100110001111010",
            data_re_out => mul_re_out(381),
            data_im_out => mul_im_out(381)
        );

 
    UMUL_382 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(382),
            data_im_in => first_stage_im_out(382),
            re_multiplicator => "0010010100101100", --- 0.580810546875 + j-0.814025878906
            im_multiplicator => "1100101111100111",
            data_re_out => mul_re_out(382),
            data_im_out => mul_im_out(382)
        );

 
    UMUL_383 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(383),
            data_im_in => first_stage_im_out(383),
            re_multiplicator => "0010010001011110", --- 0.568237304688 + j-0.822875976562
            im_multiplicator => "1100101101010110",
            data_re_out => mul_re_out(383),
            data_im_out => mul_im_out(383)
        );

 
    UMUL_384 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(384),
            data_im_in => first_stage_im_out(384),
            data_re_out => mul_re_out(384),
            data_im_out => mul_im_out(384)
        );

 
    UMUL_385 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(385),
            data_im_in => first_stage_im_out(385),
            re_multiplicator => "0011111111111101", --- 0.999816894531 + j-0.0184326171875
            im_multiplicator => "1111111011010010",
            data_re_out => mul_re_out(385),
            data_im_out => mul_im_out(385)
        );

 
    UMUL_386 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(386),
            data_im_in => first_stage_im_out(386),
            re_multiplicator => "0011111111110101", --- 0.999328613281 + j-0.0368041992188
            im_multiplicator => "1111110110100101",
            data_re_out => mul_re_out(386),
            data_im_out => mul_im_out(386)
        );

 
    UMUL_387 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(387),
            data_im_in => first_stage_im_out(387),
            re_multiplicator => "0011111111100111", --- 0.998474121094 + j-0.05517578125
            im_multiplicator => "1111110001111000",
            data_re_out => mul_re_out(387),
            data_im_out => mul_im_out(387)
        );

 
    UMUL_388 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(388),
            data_im_in => first_stage_im_out(388),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(388),
            data_im_out => mul_im_out(388)
        );

 
    UMUL_389 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(389),
            data_im_in => first_stage_im_out(389),
            re_multiplicator => "0011111110111011", --- 0.995788574219 + j-0.0919189453125
            im_multiplicator => "1111101000011110",
            data_re_out => mul_re_out(389),
            data_im_out => mul_im_out(389)
        );

 
    UMUL_390 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(390),
            data_im_in => first_stage_im_out(390),
            re_multiplicator => "0011111110011100", --- 0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(390),
            data_im_out => mul_im_out(390)
        );

 
    UMUL_391 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(391),
            data_im_in => first_stage_im_out(391),
            re_multiplicator => "0011111101111000", --- 0.99169921875 + j-0.128479003906
            im_multiplicator => "1111011111000111",
            data_re_out => mul_re_out(391),
            data_im_out => mul_im_out(391)
        );

 
    UMUL_392 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(392),
            data_im_in => first_stage_im_out(392),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(392),
            data_im_out => mul_im_out(392)
        );

 
    UMUL_393 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(393),
            data_im_in => first_stage_im_out(393),
            re_multiplicator => "0011111100100000", --- 0.986328125 + j-0.164916992188
            im_multiplicator => "1111010101110010",
            data_re_out => mul_re_out(393),
            data_im_out => mul_im_out(393)
        );

 
    UMUL_394 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(394),
            data_im_in => first_stage_im_out(394),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(394),
            data_im_out => mul_im_out(394)
        );

 
    UMUL_395 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(395),
            data_im_in => first_stage_im_out(395),
            re_multiplicator => "0011111010110001", --- 0.979553222656 + j-0.201110839844
            im_multiplicator => "1111001100100001",
            data_re_out => mul_re_out(395),
            data_im_out => mul_im_out(395)
        );

 
    UMUL_396 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(396),
            data_im_in => first_stage_im_out(396),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(396),
            data_im_out => mul_im_out(396)
        );

 
    UMUL_397 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(397),
            data_im_in => first_stage_im_out(397),
            re_multiplicator => "0011111000101101", --- 0.971496582031 + j-0.236999511719
            im_multiplicator => "1111000011010101",
            data_re_out => mul_re_out(397),
            data_im_out => mul_im_out(397)
        );

 
    UMUL_398 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(398),
            data_im_in => first_stage_im_out(398),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(398),
            data_im_out => mul_im_out(398)
        );

 
    UMUL_399 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(399),
            data_im_in => first_stage_im_out(399),
            re_multiplicator => "0011110110010011", --- 0.962097167969 + j-0.272644042969
            im_multiplicator => "1110111010001101",
            data_re_out => mul_re_out(399),
            data_im_out => mul_im_out(399)
        );

 
    UMUL_400 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(400),
            data_im_in => first_stage_im_out(400),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(400),
            data_im_out => mul_im_out(400)
        );

 
    UMUL_401 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(401),
            data_im_in => first_stage_im_out(401),
            re_multiplicator => "0011110011100100", --- 0.951416015625 + j-0.307861328125
            im_multiplicator => "1110110001001100",
            data_re_out => mul_re_out(401),
            data_im_out => mul_im_out(401)
        );

 
    UMUL_402 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(402),
            data_im_in => first_stage_im_out(402),
            re_multiplicator => "0011110010000101", --- 0.945617675781 + j-0.325317382812
            im_multiplicator => "1110101100101110",
            data_re_out => mul_re_out(402),
            data_im_out => mul_im_out(402)
        );

 
    UMUL_403 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(403),
            data_im_in => first_stage_im_out(403),
            re_multiplicator => "0011110000100000", --- 0.939453125 + j-0.342651367188
            im_multiplicator => "1110101000010010",
            data_re_out => mul_re_out(403),
            data_im_out => mul_im_out(403)
        );

 
    UMUL_404 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(404),
            data_im_in => first_stage_im_out(404),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(404),
            data_im_out => mul_im_out(404)
        );

 
    UMUL_405 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(405),
            data_im_in => first_stage_im_out(405),
            re_multiplicator => "0011101101000111", --- 0.926208496094 + j-0.377014160156
            im_multiplicator => "1110011111011111",
            data_re_out => mul_re_out(405),
            data_im_out => mul_im_out(405)
        );

 
    UMUL_406 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(406),
            data_im_in => first_stage_im_out(406),
            re_multiplicator => "0011101011010011", --- 0.919128417969 + j-0.393981933594
            im_multiplicator => "1110011011001001",
            data_re_out => mul_re_out(406),
            data_im_out => mul_im_out(406)
        );

 
    UMUL_407 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(407),
            data_im_in => first_stage_im_out(407),
            re_multiplicator => "0011101001011001", --- 0.911682128906 + j-0.410827636719
            im_multiplicator => "1110010110110101",
            data_re_out => mul_re_out(407),
            data_im_out => mul_im_out(407)
        );

 
    UMUL_408 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(408),
            data_im_in => first_stage_im_out(408),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(408),
            data_im_out => mul_im_out(408)
        );

 
    UMUL_409 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(409),
            data_im_in => first_stage_im_out(409),
            re_multiplicator => "0011100101011000", --- 0.89599609375 + j-0.444091796875
            im_multiplicator => "1110001110010100",
            data_re_out => mul_re_out(409),
            data_im_out => mul_im_out(409)
        );

 
    UMUL_410 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(410),
            data_im_in => first_stage_im_out(410),
            re_multiplicator => "0011100011001111", --- 0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(410),
            data_im_out => mul_im_out(410)
        );

 
    UMUL_411 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(411),
            data_im_in => first_stage_im_out(411),
            re_multiplicator => "0011100001000010", --- 0.879028320312 + j-0.476806640625
            im_multiplicator => "1110000101111100",
            data_re_out => mul_re_out(411),
            data_im_out => mul_im_out(411)
        );

 
    UMUL_412 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(412),
            data_im_in => first_stage_im_out(412),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(412),
            data_im_out => mul_im_out(412)
        );

 
    UMUL_413 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(413),
            data_im_in => first_stage_im_out(413),
            re_multiplicator => "0011011100011000", --- 0.86083984375 + j-0.508850097656
            im_multiplicator => "1101111101101111",
            data_re_out => mul_re_out(413),
            data_im_out => mul_im_out(413)
        );

 
    UMUL_414 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(414),
            data_im_in => first_stage_im_out(414),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(414),
            data_im_out => mul_im_out(414)
        );

 
    UMUL_415 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(415),
            data_im_in => first_stage_im_out(415),
            re_multiplicator => "0011010111011100", --- 0.841552734375 + j-0.540161132812
            im_multiplicator => "1101110101101110",
            data_re_out => mul_re_out(415),
            data_im_out => mul_im_out(415)
        );

 
    UMUL_416 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(416),
            data_im_in => first_stage_im_out(416),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(416),
            data_im_out => mul_im_out(416)
        );

 
    UMUL_417 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(417),
            data_im_in => first_stage_im_out(417),
            re_multiplicator => "0011010010001101", --- 0.821105957031 + j-0.57080078125
            im_multiplicator => "1101101101111000",
            data_re_out => mul_re_out(417),
            data_im_out => mul_im_out(417)
        );

 
    UMUL_418 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(418),
            data_im_in => first_stage_im_out(418),
            re_multiplicator => "0011001111011111", --- 0.810485839844 + j-0.585815429688
            im_multiplicator => "1101101010000010",
            data_re_out => mul_re_out(418),
            data_im_out => mul_im_out(418)
        );

 
    UMUL_419 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(419),
            data_im_in => first_stage_im_out(419),
            re_multiplicator => "0011001100101100", --- 0.799560546875 + j-0.600646972656
            im_multiplicator => "1101100110001111",
            data_re_out => mul_re_out(419),
            data_im_out => mul_im_out(419)
        );

 
    UMUL_420 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(420),
            data_im_in => first_stage_im_out(420),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(420),
            data_im_out => mul_im_out(420)
        );

 
    UMUL_421 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(421),
            data_im_in => first_stage_im_out(421),
            re_multiplicator => "0011000110111001", --- 0.776916503906 + j-0.629638671875
            im_multiplicator => "1101011110110100",
            data_re_out => mul_re_out(421),
            data_im_out => mul_im_out(421)
        );

 
    UMUL_422 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(422),
            data_im_in => first_stage_im_out(422),
            re_multiplicator => "0011000011111001", --- 0.765197753906 + j-0.643859863281
            im_multiplicator => "1101011011001011",
            data_re_out => mul_re_out(422),
            data_im_out => mul_im_out(422)
        );

 
    UMUL_423 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(423),
            data_im_in => first_stage_im_out(423),
            re_multiplicator => "0011000000110100", --- 0.753173828125 + j-0.657836914062
            im_multiplicator => "1101010111100110",
            data_re_out => mul_re_out(423),
            data_im_out => mul_im_out(423)
        );

 
    UMUL_424 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(424),
            data_im_in => first_stage_im_out(424),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(424),
            data_im_out => mul_im_out(424)
        );

 
    UMUL_425 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(425),
            data_im_in => first_stage_im_out(425),
            re_multiplicator => "0010111010011111", --- 0.728454589844 + j-0.68505859375
            im_multiplicator => "1101010000101000",
            data_re_out => mul_re_out(425),
            data_im_out => mul_im_out(425)
        );

 
    UMUL_426 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(426),
            data_im_in => first_stage_im_out(426),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(426),
            data_im_out => mul_im_out(426)
        );

 
    UMUL_427 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(427),
            data_im_in => first_stage_im_out(427),
            re_multiplicator => "0010110011111010", --- 0.702758789062 + j-0.71142578125
            im_multiplicator => "1101001001111000",
            data_re_out => mul_re_out(427),
            data_im_out => mul_im_out(427)
        );

 
    UMUL_428 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(428),
            data_im_in => first_stage_im_out(428),
            re_multiplicator => "0010110000100001", --- 0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(428),
            data_im_out => mul_im_out(428)
        );

 
    UMUL_429 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(429),
            data_im_in => first_stage_im_out(429),
            re_multiplicator => "0010101101000101", --- 0.676086425781 + j-0.73681640625
            im_multiplicator => "1101000011011000",
            data_re_out => mul_re_out(429),
            data_im_out => mul_im_out(429)
        );

 
    UMUL_430 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(430),
            data_im_in => first_stage_im_out(430),
            re_multiplicator => "0010101001100101", --- 0.662414550781 + j-0.749145507812
            im_multiplicator => "1101000000001110",
            data_re_out => mul_re_out(430),
            data_im_out => mul_im_out(430)
        );

 
    UMUL_431 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(431),
            data_im_in => first_stage_im_out(431),
            re_multiplicator => "0010100110000001", --- 0.648498535156 + j-0.76123046875
            im_multiplicator => "1100111101001000",
            data_re_out => mul_re_out(431),
            data_im_out => mul_im_out(431)
        );

 
    UMUL_432 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(432),
            data_im_in => first_stage_im_out(432),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(432),
            data_im_out => mul_im_out(432)
        );

 
    UMUL_433 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(433),
            data_im_in => first_stage_im_out(433),
            re_multiplicator => "0010011110101111", --- 0.620056152344 + j-0.784545898438
            im_multiplicator => "1100110111001010",
            data_re_out => mul_re_out(433),
            data_im_out => mul_im_out(433)
        );

 
    UMUL_434 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(434),
            data_im_in => first_stage_im_out(434),
            re_multiplicator => "0010011011000001", --- 0.605529785156 + j-0.795837402344
            im_multiplicator => "1100110100010001",
            data_re_out => mul_re_out(434),
            data_im_out => mul_im_out(434)
        );

 
    UMUL_435 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(435),
            data_im_in => first_stage_im_out(435),
            re_multiplicator => "0010010111001111", --- 0.590759277344 + j-0.806823730469
            im_multiplicator => "1100110001011101",
            data_re_out => mul_re_out(435),
            data_im_out => mul_im_out(435)
        );

 
    UMUL_436 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(436),
            data_im_in => first_stage_im_out(436),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j-0.817565917969
            im_multiplicator => "1100101110101101",
            data_re_out => mul_re_out(436),
            data_im_out => mul_im_out(436)
        );

 
    UMUL_437 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(437),
            data_im_in => first_stage_im_out(437),
            re_multiplicator => "0010001111100010", --- 0.560668945312 + j-0.828063964844
            im_multiplicator => "1100101100000001",
            data_re_out => mul_re_out(437),
            data_im_out => mul_im_out(437)
        );

 
    UMUL_438 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(438),
            data_im_in => first_stage_im_out(438),
            re_multiplicator => "0010001011100111", --- 0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(438),
            data_im_out => mul_im_out(438)
        );

 
    UMUL_439 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(439),
            data_im_in => first_stage_im_out(439),
            re_multiplicator => "0010000111101000", --- 0.52978515625 + j-0.84814453125
            im_multiplicator => "1100100110111000",
            data_re_out => mul_re_out(439),
            data_im_out => mul_im_out(439)
        );

 
    UMUL_440 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(440),
            data_im_in => first_stage_im_out(440),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(440),
            data_im_out => mul_im_out(440)
        );

 
    UMUL_441 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(441),
            data_im_in => first_stage_im_out(441),
            re_multiplicator => "0001111111100011", --- 0.498229980469 + j-0.867065429688
            im_multiplicator => "1100100010000010",
            data_re_out => mul_re_out(441),
            data_im_out => mul_im_out(441)
        );

 
    UMUL_442 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(442),
            data_im_in => first_stage_im_out(442),
            re_multiplicator => "0001111011011100", --- 0.482177734375 + j-0.876098632812
            im_multiplicator => "1100011111101110",
            data_re_out => mul_re_out(442),
            data_im_out => mul_im_out(442)
        );

 
    UMUL_443 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(443),
            data_im_in => first_stage_im_out(443),
            re_multiplicator => "0001110111010011", --- 0.466003417969 + j-0.884826660156
            im_multiplicator => "1100011101011111",
            data_re_out => mul_re_out(443),
            data_im_out => mul_im_out(443)
        );

 
    UMUL_444 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(444),
            data_im_in => first_stage_im_out(444),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(444),
            data_im_out => mul_im_out(444)
        );

 
    UMUL_445 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(445),
            data_im_in => first_stage_im_out(445),
            re_multiplicator => "0001101110111000", --- 0.43310546875 + j-0.9013671875
            im_multiplicator => "1100011001010000",
            data_re_out => mul_re_out(445),
            data_im_out => mul_im_out(445)
        );

 
    UMUL_446 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(446),
            data_im_in => first_stage_im_out(446),
            re_multiplicator => "0001101010100111", --- 0.416442871094 + j-0.9091796875
            im_multiplicator => "1100010111010000",
            data_re_out => mul_re_out(446),
            data_im_out => mul_im_out(446)
        );

 
    UMUL_447 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(447),
            data_im_in => first_stage_im_out(447),
            re_multiplicator => "0001100110010011", --- 0.399597167969 + j-0.916687011719
            im_multiplicator => "1100010101010101",
            data_re_out => mul_re_out(447),
            data_im_out => mul_im_out(447)
        );

 
    UMUL_448 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(448),
            data_im_in => first_stage_im_out(448),
            data_re_out => mul_re_out(448),
            data_im_out => mul_im_out(448)
        );

 
    UMUL_449 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(449),
            data_im_in => first_stage_im_out(449),
            re_multiplicator => "0011111111111100", --- 0.999755859375 + j-0.021484375
            im_multiplicator => "1111111010100000",
            data_re_out => mul_re_out(449),
            data_im_out => mul_im_out(449)
        );

 
    UMUL_450 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(450),
            data_im_in => first_stage_im_out(450),
            re_multiplicator => "0011111111110001", --- 0.999084472656 + j-0.04296875
            im_multiplicator => "1111110101000000",
            data_re_out => mul_re_out(450),
            data_im_out => mul_im_out(450)
        );

 
    UMUL_451 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(451),
            data_im_in => first_stage_im_out(451),
            re_multiplicator => "0011111111011110", --- 0.997924804688 + j-0.0643920898438
            im_multiplicator => "1111101111100001",
            data_re_out => mul_re_out(451),
            data_im_out => mul_im_out(451)
        );

 
    UMUL_452 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(452),
            data_im_in => first_stage_im_out(452),
            re_multiplicator => "0011111111000100", --- 0.996337890625 + j-0.0858154296875
            im_multiplicator => "1111101010000010",
            data_re_out => mul_re_out(452),
            data_im_out => mul_im_out(452)
        );

 
    UMUL_453 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(453),
            data_im_in => first_stage_im_out(453),
            re_multiplicator => "0011111110100010", --- 0.994262695312 + j-0.107177734375
            im_multiplicator => "1111100100100100",
            data_re_out => mul_re_out(453),
            data_im_out => mul_im_out(453)
        );

 
    UMUL_454 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(454),
            data_im_in => first_stage_im_out(454),
            re_multiplicator => "0011111101111000", --- 0.99169921875 + j-0.128479003906
            im_multiplicator => "1111011111000111",
            data_re_out => mul_re_out(454),
            data_im_out => mul_im_out(454)
        );

 
    UMUL_455 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(455),
            data_im_in => first_stage_im_out(455),
            re_multiplicator => "0011111101000111", --- 0.988708496094 + j-0.149780273438
            im_multiplicator => "1111011001101010",
            data_re_out => mul_re_out(455),
            data_im_out => mul_im_out(455)
        );

 
    UMUL_456 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(456),
            data_im_in => first_stage_im_out(456),
            re_multiplicator => "0011111100001111", --- 0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(456),
            data_im_out => mul_im_out(456)
        );

 
    UMUL_457 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(457),
            data_im_in => first_stage_im_out(457),
            re_multiplicator => "0011111011001111", --- 0.981384277344 + j-0.192077636719
            im_multiplicator => "1111001110110101",
            data_re_out => mul_re_out(457),
            data_im_out => mul_im_out(457)
        );

 
    UMUL_458 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(458),
            data_im_in => first_stage_im_out(458),
            re_multiplicator => "0011111010001000", --- 0.97705078125 + j-0.213134765625
            im_multiplicator => "1111001001011100",
            data_re_out => mul_re_out(458),
            data_im_out => mul_im_out(458)
        );

 
    UMUL_459 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(459),
            data_im_in => first_stage_im_out(459),
            re_multiplicator => "0011111000111001", --- 0.972229003906 + j-0.234069824219
            im_multiplicator => "1111000100000101",
            data_re_out => mul_re_out(459),
            data_im_out => mul_im_out(459)
        );

 
    UMUL_460 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(460),
            data_im_in => first_stage_im_out(460),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(460),
            data_im_out => mul_im_out(460)
        );

 
    UMUL_461 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(461),
            data_im_in => first_stage_im_out(461),
            re_multiplicator => "0011110110000110", --- 0.961303710938 + j-0.275573730469
            im_multiplicator => "1110111001011101",
            data_re_out => mul_re_out(461),
            data_im_out => mul_im_out(461)
        );

 
    UMUL_462 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(462),
            data_im_in => first_stage_im_out(462),
            re_multiplicator => "0011110100100001", --- 0.955139160156 + j-0.296142578125
            im_multiplicator => "1110110100001100",
            data_re_out => mul_re_out(462),
            data_im_out => mul_im_out(462)
        );

 
    UMUL_463 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(463),
            data_im_in => first_stage_im_out(463),
            re_multiplicator => "0011110010110101", --- 0.948547363281 + j-0.316589355469
            im_multiplicator => "1110101110111101",
            data_re_out => mul_re_out(463),
            data_im_out => mul_im_out(463)
        );

 
    UMUL_464 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(464),
            data_im_in => first_stage_im_out(464),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(464),
            data_im_out => mul_im_out(464)
        );

 
    UMUL_465 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(465),
            data_im_in => first_stage_im_out(465),
            re_multiplicator => "0011101111001000", --- 0.93408203125 + j-0.357055664062
            im_multiplicator => "1110100100100110",
            data_re_out => mul_re_out(465),
            data_im_out => mul_im_out(465)
        );

 
    UMUL_466 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(466),
            data_im_in => first_stage_im_out(466),
            re_multiplicator => "0011101101000111", --- 0.926208496094 + j-0.377014160156
            im_multiplicator => "1110011111011111",
            data_re_out => mul_re_out(466),
            data_im_out => mul_im_out(466)
        );

 
    UMUL_467 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(467),
            data_im_in => first_stage_im_out(467),
            re_multiplicator => "0011101010111111", --- 0.917907714844 + j-0.396789550781
            im_multiplicator => "1110011010011011",
            data_re_out => mul_re_out(467),
            data_im_out => mul_im_out(467)
        );

 
    UMUL_468 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(468),
            data_im_in => first_stage_im_out(468),
            re_multiplicator => "0011101000110000", --- 0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(468),
            data_im_out => mul_im_out(468)
        );

 
    UMUL_469 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(469),
            data_im_in => first_stage_im_out(469),
            re_multiplicator => "0011100110011010", --- 0.900024414062 + j-0.435852050781
            im_multiplicator => "1110010000011011",
            data_re_out => mul_re_out(469),
            data_im_out => mul_im_out(469)
        );

 
    UMUL_470 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(470),
            data_im_in => first_stage_im_out(470),
            re_multiplicator => "0011100011111101", --- 0.890441894531 + j-0.455078125
            im_multiplicator => "1110001011100000",
            data_re_out => mul_re_out(470),
            data_im_out => mul_im_out(470)
        );

 
    UMUL_471 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(471),
            data_im_in => first_stage_im_out(471),
            re_multiplicator => "0011100001011010", --- 0.880493164062 + j-0.47412109375
            im_multiplicator => "1110000110101000",
            data_re_out => mul_re_out(471),
            data_im_out => mul_im_out(471)
        );

 
    UMUL_472 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(472),
            data_im_in => first_stage_im_out(472),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(472),
            data_im_out => mul_im_out(472)
        );

 
    UMUL_473 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(473),
            data_im_in => first_stage_im_out(473),
            re_multiplicator => "0011011011111111", --- 0.859313964844 + j-0.511474609375
            im_multiplicator => "1101111101000100",
            data_re_out => mul_re_out(473),
            data_im_out => mul_im_out(473)
        );

 
    UMUL_474 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(474),
            data_im_in => first_stage_im_out(474),
            re_multiplicator => "0011011001001000", --- 0.84814453125 + j-0.52978515625
            im_multiplicator => "1101111000011000",
            data_re_out => mul_re_out(474),
            data_im_out => mul_im_out(474)
        );

 
    UMUL_475 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(475),
            data_im_in => first_stage_im_out(475),
            re_multiplicator => "0011010110001010", --- 0.836547851562 + j-0.547912597656
            im_multiplicator => "1101110011101111",
            data_re_out => mul_re_out(475),
            data_im_out => mul_im_out(475)
        );

 
    UMUL_476 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(476),
            data_im_in => first_stage_im_out(476),
            re_multiplicator => "0011010011000110", --- 0.824584960938 + j-0.565734863281
            im_multiplicator => "1101101111001011",
            data_re_out => mul_re_out(476),
            data_im_out => mul_im_out(476)
        );

 
    UMUL_477 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(477),
            data_im_in => first_stage_im_out(477),
            re_multiplicator => "0011001111111100", --- 0.812255859375 + j-0.583312988281
            im_multiplicator => "1101101010101011",
            data_re_out => mul_re_out(477),
            data_im_out => mul_im_out(477)
        );

 
    UMUL_478 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(478),
            data_im_in => first_stage_im_out(478),
            re_multiplicator => "0011001100101100", --- 0.799560546875 + j-0.600646972656
            im_multiplicator => "1101100110001111",
            data_re_out => mul_re_out(478),
            data_im_out => mul_im_out(478)
        );

 
    UMUL_479 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(479),
            data_im_in => first_stage_im_out(479),
            re_multiplicator => "0011001001010101", --- 0.786437988281 + j-0.61767578125
            im_multiplicator => "1101100001111000",
            data_re_out => mul_re_out(479),
            data_im_out => mul_im_out(479)
        );

 
    UMUL_480 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(480),
            data_im_in => first_stage_im_out(480),
            re_multiplicator => "0011000101111001", --- 0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(480),
            data_im_out => mul_im_out(480)
        );

 
    UMUL_481 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(481),
            data_im_in => first_stage_im_out(481),
            re_multiplicator => "0011000010010111", --- 0.759216308594 + j-0.650817871094
            im_multiplicator => "1101011001011001",
            data_re_out => mul_re_out(481),
            data_im_out => mul_im_out(481)
        );

 
    UMUL_482 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(482),
            data_im_in => first_stage_im_out(482),
            re_multiplicator => "0010111110101111", --- 0.745056152344 + j-0.6669921875
            im_multiplicator => "1101010101010000",
            data_re_out => mul_re_out(482),
            data_im_out => mul_im_out(482)
        );

 
    UMUL_483 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(483),
            data_im_in => first_stage_im_out(483),
            re_multiplicator => "0010111011000010", --- 0.730590820312 + j-0.682861328125
            im_multiplicator => "1101010001001100",
            data_re_out => mul_re_out(483),
            data_im_out => mul_im_out(483)
        );

 
    UMUL_484 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(484),
            data_im_in => first_stage_im_out(484),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(484),
            data_im_out => mul_im_out(484)
        );

 
    UMUL_485 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(485),
            data_im_in => first_stage_im_out(485),
            re_multiplicator => "0010110011010110", --- 0.700561523438 + j-0.713562011719
            im_multiplicator => "1101001001010101",
            data_re_out => mul_re_out(485),
            data_im_out => mul_im_out(485)
        );

 
    UMUL_486 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(486),
            data_im_in => first_stage_im_out(486),
            re_multiplicator => "0010101111011000", --- 0.68505859375 + j-0.728454589844
            im_multiplicator => "1101000101100001",
            data_re_out => mul_re_out(486),
            data_im_out => mul_im_out(486)
        );

 
    UMUL_487 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(487),
            data_im_in => first_stage_im_out(487),
            re_multiplicator => "0010101011010110", --- 0.669311523438 + j-0.742980957031
            im_multiplicator => "1101000001110011",
            data_re_out => mul_re_out(487),
            data_im_out => mul_im_out(487)
        );

 
    UMUL_488 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(488),
            data_im_in => first_stage_im_out(488),
            re_multiplicator => "0010100111001110", --- 0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(488),
            data_im_out => mul_im_out(488)
        );

 
    UMUL_489 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(489),
            data_im_in => first_stage_im_out(489),
            re_multiplicator => "0010100011000001", --- 0.636779785156 + j-0.771057128906
            im_multiplicator => "1100111010100111",
            data_re_out => mul_re_out(489),
            data_im_out => mul_im_out(489)
        );

 
    UMUL_490 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(490),
            data_im_in => first_stage_im_out(490),
            re_multiplicator => "0010011110101111", --- 0.620056152344 + j-0.784545898438
            im_multiplicator => "1100110111001010",
            data_re_out => mul_re_out(490),
            data_im_out => mul_im_out(490)
        );

 
    UMUL_491 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(491),
            data_im_in => first_stage_im_out(491),
            re_multiplicator => "0010011010011001", --- 0.603088378906 + j-0.797668457031
            im_multiplicator => "1100110011110011",
            data_re_out => mul_re_out(491),
            data_im_out => mul_im_out(491)
        );

 
    UMUL_492 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(492),
            data_im_in => first_stage_im_out(492),
            re_multiplicator => "0010010101111110", --- 0.585815429688 + j-0.810485839844
            im_multiplicator => "1100110000100001",
            data_re_out => mul_re_out(492),
            data_im_out => mul_im_out(492)
        );

 
    UMUL_493 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(493),
            data_im_in => first_stage_im_out(493),
            re_multiplicator => "0010010001011110", --- 0.568237304688 + j-0.822875976562
            im_multiplicator => "1100101101010110",
            data_re_out => mul_re_out(493),
            data_im_out => mul_im_out(493)
        );

 
    UMUL_494 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(494),
            data_im_in => first_stage_im_out(494),
            re_multiplicator => "0010001100111011", --- 0.550476074219 + j-0.834838867188
            im_multiplicator => "1100101010010010",
            data_re_out => mul_re_out(494),
            data_im_out => mul_im_out(494)
        );

 
    UMUL_495 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(495),
            data_im_in => first_stage_im_out(495),
            re_multiplicator => "0010001000010011", --- 0.532409667969 + j-0.846496582031
            im_multiplicator => "1100100111010011",
            data_re_out => mul_re_out(495),
            data_im_out => mul_im_out(495)
        );

 
    UMUL_496 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(496),
            data_im_in => first_stage_im_out(496),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(496),
            data_im_out => mul_im_out(496)
        );

 
    UMUL_497 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(497),
            data_im_in => first_stage_im_out(497),
            re_multiplicator => "0001111110110111", --- 0.495544433594 + j-0.868591308594
            im_multiplicator => "1100100001101001",
            data_re_out => mul_re_out(497),
            data_im_out => mul_im_out(497)
        );

 
    UMUL_498 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(498),
            data_im_in => first_stage_im_out(498),
            re_multiplicator => "0001111010000100", --- 0.476806640625 + j-0.879028320312
            im_multiplicator => "1100011110111110",
            data_re_out => mul_re_out(498),
            data_im_out => mul_im_out(498)
        );

 
    UMUL_499 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(499),
            data_im_in => first_stage_im_out(499),
            re_multiplicator => "0001110101001101", --- 0.457824707031 + j-0.889038085938
            im_multiplicator => "1100011100011010",
            data_re_out => mul_re_out(499),
            data_im_out => mul_im_out(499)
        );

 
    UMUL_500 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(500),
            data_im_in => first_stage_im_out(500),
            re_multiplicator => "0001110000010010", --- 0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(500),
            data_im_out => mul_im_out(500)
        );

 
    UMUL_501 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(501),
            data_im_in => first_stage_im_out(501),
            re_multiplicator => "0001101011010100", --- 0.419189453125 + j-0.907897949219
            im_multiplicator => "1100010111100101",
            data_re_out => mul_re_out(501),
            data_im_out => mul_im_out(501)
        );

 
    UMUL_502 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(502),
            data_im_in => first_stage_im_out(502),
            re_multiplicator => "0001100110010011", --- 0.399597167969 + j-0.916687011719
            im_multiplicator => "1100010101010101",
            data_re_out => mul_re_out(502),
            data_im_out => mul_im_out(502)
        );

 
    UMUL_503 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(503),
            data_im_in => first_stage_im_out(503),
            re_multiplicator => "0001100001001111", --- 0.379821777344 + j-0.925048828125
            im_multiplicator => "1100010011001100",
            data_re_out => mul_re_out(503),
            data_im_out => mul_im_out(503)
        );

 
    UMUL_504 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(504),
            data_im_in => first_stage_im_out(504),
            re_multiplicator => "0001011100001001", --- 0.359924316406 + j-0.932983398438
            im_multiplicator => "1100010001001010",
            data_re_out => mul_re_out(504),
            data_im_out => mul_im_out(504)
        );

 
    UMUL_505 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(505),
            data_im_in => first_stage_im_out(505),
            re_multiplicator => "0001010110111111", --- 0.339782714844 + j-0.940490722656
            im_multiplicator => "1100001111001111",
            data_re_out => mul_re_out(505),
            data_im_out => mul_im_out(505)
        );

 
    UMUL_506 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(506),
            data_im_in => first_stage_im_out(506),
            re_multiplicator => "0001010001110011", --- 0.319519042969 + j-0.947570800781
            im_multiplicator => "1100001101011011",
            data_re_out => mul_re_out(506),
            data_im_out => mul_im_out(506)
        );

 
    UMUL_507 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(507),
            data_im_in => first_stage_im_out(507),
            re_multiplicator => "0001001100100100", --- 0.299072265625 + j-0.954223632812
            im_multiplicator => "1100001011101110",
            data_re_out => mul_re_out(507),
            data_im_out => mul_im_out(507)
        );

 
    UMUL_508 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(508),
            data_im_in => first_stage_im_out(508),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(508),
            data_im_out => mul_im_out(508)
        );

 
    UMUL_509 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(509),
            data_im_in => first_stage_im_out(509),
            re_multiplicator => "0001000010000000", --- 0.2578125 + j-0.966186523438
            im_multiplicator => "1100001000101010",
            data_re_out => mul_re_out(509),
            data_im_out => mul_im_out(509)
        );

 
    UMUL_510 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(510),
            data_im_in => first_stage_im_out(510),
            re_multiplicator => "0000111100101011", --- 0.236999511719 + j-0.971496582031
            im_multiplicator => "1100000111010011",
            data_re_out => mul_re_out(510),
            data_im_out => mul_im_out(510)
        );

 
    UMUL_511 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(511),
            data_im_in => first_stage_im_out(511),
            re_multiplicator => "0000110111010101", --- 0.216125488281 + j-0.976379394531
            im_multiplicator => "1100000110000011",
            data_re_out => mul_re_out(511),
            data_im_out => mul_im_out(511)
        );

 
    UMUL_512 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(512),
            data_im_in => first_stage_im_out(512),
            data_re_out => mul_re_out(512),
            data_im_out => mul_im_out(512)
        );

 
    UMUL_513 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(513),
            data_im_in => first_stage_im_out(513),
            re_multiplicator => "0011111111111011", --- 0.999694824219 + j-0.0245361328125
            im_multiplicator => "1111111001101110",
            data_re_out => mul_re_out(513),
            data_im_out => mul_im_out(513)
        );

 
    UMUL_514 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(514),
            data_im_in => first_stage_im_out(514),
            re_multiplicator => "0011111111101100", --- 0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(514),
            data_im_out => mul_im_out(514)
        );

 
    UMUL_515 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(515),
            data_im_in => first_stage_im_out(515),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(515),
            data_im_out => mul_im_out(515)
        );

 
    UMUL_516 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(516),
            data_im_in => first_stage_im_out(516),
            re_multiplicator => "0011111110110001", --- 0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(516),
            data_im_out => mul_im_out(516)
        );

 
    UMUL_517 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(517),
            data_im_in => first_stage_im_out(517),
            re_multiplicator => "0011111110000101", --- 0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(517),
            data_im_out => mul_im_out(517)
        );

 
    UMUL_518 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(518),
            data_im_in => first_stage_im_out(518),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(518),
            data_im_out => mul_im_out(518)
        );

 
    UMUL_519 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(519),
            data_im_in => first_stage_im_out(519),
            re_multiplicator => "0011111100001111", --- 0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(519),
            data_im_out => mul_im_out(519)
        );

 
    UMUL_520 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(520),
            data_im_in => first_stage_im_out(520),
            re_multiplicator => "0011111011000101", --- 0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(520),
            data_im_out => mul_im_out(520)
        );

 
    UMUL_521 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(521),
            data_im_in => first_stage_im_out(521),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(521),
            data_im_out => mul_im_out(521)
        );

 
    UMUL_522 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(522),
            data_im_in => first_stage_im_out(522),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(522),
            data_im_out => mul_im_out(522)
        );

 
    UMUL_523 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(523),
            data_im_in => first_stage_im_out(523),
            re_multiplicator => "0011110110101111", --- 0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(523),
            data_im_out => mul_im_out(523)
        );

 
    UMUL_524 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(524),
            data_im_in => first_stage_im_out(524),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(524),
            data_im_out => mul_im_out(524)
        );

 
    UMUL_525 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(525),
            data_im_in => first_stage_im_out(525),
            re_multiplicator => "0011110011000101", --- 0.949523925781 + j-0.313659667969
            im_multiplicator => "1110101111101101",
            data_re_out => mul_re_out(525),
            data_im_out => mul_im_out(525)
        );

 
    UMUL_526 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(526),
            data_im_in => first_stage_im_out(526),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(526),
            data_im_out => mul_im_out(526)
        );

 
    UMUL_527 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(527),
            data_im_in => first_stage_im_out(527),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(527),
            data_im_out => mul_im_out(527)
        );

 
    UMUL_528 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(528),
            data_im_in => first_stage_im_out(528),
            re_multiplicator => "0011101100100001", --- 0.923889160156 + j-0.382690429688
            im_multiplicator => "1110011110000010",
            data_re_out => mul_re_out(528),
            data_im_out => mul_im_out(528)
        );

 
    UMUL_529 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(529),
            data_im_in => first_stage_im_out(529),
            re_multiplicator => "0011101010000010", --- 0.914184570312 + j-0.405212402344
            im_multiplicator => "1110011000010001",
            data_re_out => mul_re_out(529),
            data_im_out => mul_im_out(529)
        );

 
    UMUL_530 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(530),
            data_im_in => first_stage_im_out(530),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(530),
            data_im_out => mul_im_out(530)
        );

 
    UMUL_531 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(531),
            data_im_in => first_stage_im_out(531),
            re_multiplicator => "0011100100101011", --- 0.893249511719 + j-0.449584960938
            im_multiplicator => "1110001100111010",
            data_re_out => mul_re_out(531),
            data_im_out => mul_im_out(531)
        );

 
    UMUL_532 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(532),
            data_im_in => first_stage_im_out(532),
            re_multiplicator => "0011100001110001", --- 0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(532),
            data_im_out => mul_im_out(532)
        );

 
    UMUL_533 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(533),
            data_im_in => first_stage_im_out(533),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(533),
            data_im_out => mul_im_out(533)
        );

 
    UMUL_534 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(534),
            data_im_in => first_stage_im_out(534),
            re_multiplicator => "0011011011100101", --- 0.857727050781 + j-0.514099121094
            im_multiplicator => "1101111100011001",
            data_re_out => mul_re_out(534),
            data_im_out => mul_im_out(534)
        );

 
    UMUL_535 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(535),
            data_im_in => first_stage_im_out(535),
            re_multiplicator => "0011011000010010", --- 0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(535),
            data_im_out => mul_im_out(535)
        );

 
    UMUL_536 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(536),
            data_im_in => first_stage_im_out(536),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(536),
            data_im_out => mul_im_out(536)
        );

 
    UMUL_537 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(537),
            data_im_in => first_stage_im_out(537),
            re_multiplicator => "0011010001010011", --- 0.817565917969 + j-0.575805664062
            im_multiplicator => "1101101100100110",
            data_re_out => mul_re_out(537),
            data_im_out => mul_im_out(537)
        );

 
    UMUL_538 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(538),
            data_im_in => first_stage_im_out(538),
            re_multiplicator => "0011001101101000", --- 0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(538),
            data_im_out => mul_im_out(538)
        );

 
    UMUL_539 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(539),
            data_im_in => first_stage_im_out(539),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(539),
            data_im_out => mul_im_out(539)
        );

 
    UMUL_540 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(540),
            data_im_in => first_stage_im_out(540),
            re_multiplicator => "0011000101111001", --- 0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(540),
            data_im_out => mul_im_out(540)
        );

 
    UMUL_541 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(541),
            data_im_in => first_stage_im_out(541),
            re_multiplicator => "0011000001110110", --- 0.757202148438 + j-0.653198242188
            im_multiplicator => "1101011000110010",
            data_re_out => mul_re_out(541),
            data_im_out => mul_im_out(541)
        );

 
    UMUL_542 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(542),
            data_im_in => first_stage_im_out(542),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(542),
            data_im_out => mul_im_out(542)
        );

 
    UMUL_543 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(543),
            data_im_in => first_stage_im_out(543),
            re_multiplicator => "0010111001011010", --- 0.724243164062 + j-0.689514160156
            im_multiplicator => "1101001111011111",
            data_re_out => mul_re_out(543),
            data_im_out => mul_im_out(543)
        );

 
    UMUL_544 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(544),
            data_im_in => first_stage_im_out(544),
            re_multiplicator => "0010110101000001", --- 0.707092285156 + j-0.707092285156
            im_multiplicator => "1101001010111111",
            data_re_out => mul_re_out(544),
            data_im_out => mul_im_out(544)
        );

 
    UMUL_545 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(545),
            data_im_in => first_stage_im_out(545),
            re_multiplicator => "0010110000100001", --- 0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(545),
            data_im_out => mul_im_out(545)
        );

 
    UMUL_546 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(546),
            data_im_in => first_stage_im_out(546),
            re_multiplicator => "0010101011111011", --- 0.671569824219 + j-0.740966796875
            im_multiplicator => "1101000010010100",
            data_re_out => mul_re_out(546),
            data_im_out => mul_im_out(546)
        );

 
    UMUL_547 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(547),
            data_im_in => first_stage_im_out(547),
            re_multiplicator => "0010100111001110", --- 0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(547),
            data_im_out => mul_im_out(547)
        );

 
    UMUL_548 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(548),
            data_im_in => first_stage_im_out(548),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(548),
            data_im_out => mul_im_out(548)
        );

 
    UMUL_549 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(549),
            data_im_in => first_stage_im_out(549),
            re_multiplicator => "0010011101100000", --- 0.615234375 + j-0.788330078125
            im_multiplicator => "1100110110001100",
            data_re_out => mul_re_out(549),
            data_im_out => mul_im_out(549)
        );

 
    UMUL_550 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(550),
            data_im_in => first_stage_im_out(550),
            re_multiplicator => "0010011000100000", --- 0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(550),
            data_im_out => mul_im_out(550)
        );

 
    UMUL_551 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(551),
            data_im_in => first_stage_im_out(551),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j-0.817565917969
            im_multiplicator => "1100101110101101",
            data_re_out => mul_re_out(551),
            data_im_out => mul_im_out(551)
        );

 
    UMUL_552 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(552),
            data_im_in => first_stage_im_out(552),
            re_multiplicator => "0010001110001110", --- 0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(552),
            data_im_out => mul_im_out(552)
        );

 
    UMUL_553 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(553),
            data_im_in => first_stage_im_out(553),
            re_multiplicator => "0010001000111101", --- 0.534973144531 + j-0.844848632812
            im_multiplicator => "1100100111101110",
            data_re_out => mul_re_out(553),
            data_im_out => mul_im_out(553)
        );

 
    UMUL_554 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(554),
            data_im_in => first_stage_im_out(554),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(554),
            data_im_out => mul_im_out(554)
        );

 
    UMUL_555 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(555),
            data_im_in => first_stage_im_out(555),
            re_multiplicator => "0001111110001100", --- 0.492919921875 + j-0.8701171875
            im_multiplicator => "1100100001010000",
            data_re_out => mul_re_out(555),
            data_im_out => mul_im_out(555)
        );

 
    UMUL_556 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(556),
            data_im_in => first_stage_im_out(556),
            re_multiplicator => "0001111000101011", --- 0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(556),
            data_im_out => mul_im_out(556)
        );

 
    UMUL_557 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(557),
            data_im_in => first_stage_im_out(557),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(557),
            data_im_out => mul_im_out(557)
        );

 
    UMUL_558 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(558),
            data_im_in => first_stage_im_out(558),
            re_multiplicator => "0001101101011101", --- 0.427551269531 + j-0.903991699219
            im_multiplicator => "1100011000100101",
            data_re_out => mul_re_out(558),
            data_im_out => mul_im_out(558)
        );

 
    UMUL_559 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(559),
            data_im_in => first_stage_im_out(559),
            re_multiplicator => "0001100111101111", --- 0.405212402344 + j-0.914184570312
            im_multiplicator => "1100010101111110",
            data_re_out => mul_re_out(559),
            data_im_out => mul_im_out(559)
        );

 
    UMUL_560 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(560),
            data_im_in => first_stage_im_out(560),
            re_multiplicator => "0001100001111110", --- 0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(560),
            data_im_out => mul_im_out(560)
        );

 
    UMUL_561 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(561),
            data_im_in => first_stage_im_out(561),
            re_multiplicator => "0001011100001001", --- 0.359924316406 + j-0.932983398438
            im_multiplicator => "1100010001001010",
            data_re_out => mul_re_out(561),
            data_im_out => mul_im_out(561)
        );

 
    UMUL_562 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(562),
            data_im_in => first_stage_im_out(562),
            re_multiplicator => "0001010110010000", --- 0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(562),
            data_im_out => mul_im_out(562)
        );

 
    UMUL_563 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(563),
            data_im_in => first_stage_im_out(563),
            re_multiplicator => "0001010000010011", --- 0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(563),
            data_im_out => mul_im_out(563)
        );

 
    UMUL_564 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(564),
            data_im_in => first_stage_im_out(564),
            re_multiplicator => "0001001010010100", --- 0.290283203125 + j-0.956970214844
            im_multiplicator => "1100001011000001",
            data_re_out => mul_re_out(564),
            data_im_out => mul_im_out(564)
        );

 
    UMUL_565 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(565),
            data_im_in => first_stage_im_out(565),
            re_multiplicator => "0001000100010010", --- 0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(565),
            data_im_out => mul_im_out(565)
        );

 
    UMUL_566 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(566),
            data_im_in => first_stage_im_out(566),
            re_multiplicator => "0000111110001101", --- 0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(566),
            data_im_out => mul_im_out(566)
        );

 
    UMUL_567 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(567),
            data_im_in => first_stage_im_out(567),
            re_multiplicator => "0000111000000110", --- 0.219116210938 + j-0.975708007812
            im_multiplicator => "1100000110001110",
            data_re_out => mul_re_out(567),
            data_im_out => mul_im_out(567)
        );

 
    UMUL_568 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(568),
            data_im_in => first_stage_im_out(568),
            re_multiplicator => "0000110001111100", --- 0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(568),
            data_im_out => mul_im_out(568)
        );

 
    UMUL_569 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(569),
            data_im_in => first_stage_im_out(569),
            re_multiplicator => "0000101011110001", --- 0.170959472656 + j-0.985290527344
            im_multiplicator => "1100000011110001",
            data_re_out => mul_re_out(569),
            data_im_out => mul_im_out(569)
        );

 
    UMUL_570 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(570),
            data_im_in => first_stage_im_out(570),
            re_multiplicator => "0000100101100100", --- 0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(570),
            data_im_out => mul_im_out(570)
        );

 
    UMUL_571 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(571),
            data_im_in => first_stage_im_out(571),
            re_multiplicator => "0000011111010110", --- 0.122436523438 + j-0.992492675781
            im_multiplicator => "1100000001111011",
            data_re_out => mul_re_out(571),
            data_im_out => mul_im_out(571)
        );

 
    UMUL_572 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(572),
            data_im_in => first_stage_im_out(572),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(572),
            data_im_out => mul_im_out(572)
        );

 
    UMUL_573 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(573),
            data_im_in => first_stage_im_out(573),
            re_multiplicator => "0000010010110101", --- 0.0735473632812 + j-0.997314453125
            im_multiplicator => "1100000000101100",
            data_re_out => mul_re_out(573),
            data_im_out => mul_im_out(573)
        );

 
    UMUL_574 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(574),
            data_im_in => first_stage_im_out(574),
            re_multiplicator => "0000001100100100", --- 0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(574),
            data_im_out => mul_im_out(574)
        );

 
    UMUL_575 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(575),
            data_im_in => first_stage_im_out(575),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(575),
            data_im_out => mul_im_out(575)
        );

 
    UMUL_576 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(576),
            data_im_in => first_stage_im_out(576),
            data_re_out => mul_re_out(576),
            data_im_out => mul_im_out(576)
        );

 
    UMUL_577 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(577),
            data_im_in => first_stage_im_out(577),
            re_multiplicator => "0011111111111010", --- 0.999633789062 + j-0.027587890625
            im_multiplicator => "1111111000111100",
            data_re_out => mul_re_out(577),
            data_im_out => mul_im_out(577)
        );

 
    UMUL_578 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(578),
            data_im_in => first_stage_im_out(578),
            re_multiplicator => "0011111111100111", --- 0.998474121094 + j-0.05517578125
            im_multiplicator => "1111110001111000",
            data_re_out => mul_re_out(578),
            data_im_out => mul_im_out(578)
        );

 
    UMUL_579 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(579),
            data_im_in => first_stage_im_out(579),
            re_multiplicator => "0011111111001000", --- 0.99658203125 + j-0.082763671875
            im_multiplicator => "1111101010110100",
            data_re_out => mul_re_out(579),
            data_im_out => mul_im_out(579)
        );

 
    UMUL_580 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(580),
            data_im_in => first_stage_im_out(580),
            re_multiplicator => "0011111110011100", --- 0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(580),
            data_im_out => mul_im_out(580)
        );

 
    UMUL_581 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(581),
            data_im_in => first_stage_im_out(581),
            re_multiplicator => "0011111101100100", --- 0.990478515625 + j-0.137634277344
            im_multiplicator => "1111011100110001",
            data_re_out => mul_re_out(581),
            data_im_out => mul_im_out(581)
        );

 
    UMUL_582 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(582),
            data_im_in => first_stage_im_out(582),
            re_multiplicator => "0011111100100000", --- 0.986328125 + j-0.164916992188
            im_multiplicator => "1111010101110010",
            data_re_out => mul_re_out(582),
            data_im_out => mul_im_out(582)
        );

 
    UMUL_583 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(583),
            data_im_in => first_stage_im_out(583),
            re_multiplicator => "0011111011001111", --- 0.981384277344 + j-0.192077636719
            im_multiplicator => "1111001110110101",
            data_re_out => mul_re_out(583),
            data_im_out => mul_im_out(583)
        );

 
    UMUL_584 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(584),
            data_im_in => first_stage_im_out(584),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(584),
            data_im_out => mul_im_out(584)
        );

 
    UMUL_585 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(585),
            data_im_in => first_stage_im_out(585),
            re_multiplicator => "0011111000001001", --- 0.969299316406 + j-0.245971679688
            im_multiplicator => "1111000001000010",
            data_re_out => mul_re_out(585),
            data_im_out => mul_im_out(585)
        );

 
    UMUL_586 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(586),
            data_im_in => first_stage_im_out(586),
            re_multiplicator => "0011110110010011", --- 0.962097167969 + j-0.272644042969
            im_multiplicator => "1110111010001101",
            data_re_out => mul_re_out(586),
            data_im_out => mul_im_out(586)
        );

 
    UMUL_587 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(587),
            data_im_in => first_stage_im_out(587),
            re_multiplicator => "0011110100010010", --- 0.954223632812 + j-0.299072265625
            im_multiplicator => "1110110011011100",
            data_re_out => mul_re_out(587),
            data_im_out => mul_im_out(587)
        );

 
    UMUL_588 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(588),
            data_im_in => first_stage_im_out(588),
            re_multiplicator => "0011110010000101", --- 0.945617675781 + j-0.325317382812
            im_multiplicator => "1110101100101110",
            data_re_out => mul_re_out(588),
            data_im_out => mul_im_out(588)
        );

 
    UMUL_589 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(589),
            data_im_in => first_stage_im_out(589),
            re_multiplicator => "0011101111101100", --- 0.936279296875 + j-0.351318359375
            im_multiplicator => "1110100110000100",
            data_re_out => mul_re_out(589),
            data_im_out => mul_im_out(589)
        );

 
    UMUL_590 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(590),
            data_im_in => first_stage_im_out(590),
            re_multiplicator => "0011101101000111", --- 0.926208496094 + j-0.377014160156
            im_multiplicator => "1110011111011111",
            data_re_out => mul_re_out(590),
            data_im_out => mul_im_out(590)
        );

 
    UMUL_591 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(591),
            data_im_in => first_stage_im_out(591),
            re_multiplicator => "0011101010010111", --- 0.915466308594 + j-0.402404785156
            im_multiplicator => "1110011000111111",
            data_re_out => mul_re_out(591),
            data_im_out => mul_im_out(591)
        );

 
    UMUL_592 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(592),
            data_im_in => first_stage_im_out(592),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(592),
            data_im_out => mul_im_out(592)
        );

 
    UMUL_593 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(593),
            data_im_in => first_stage_im_out(593),
            re_multiplicator => "0011100100010100", --- 0.891845703125 + j-0.452331542969
            im_multiplicator => "1110001100001101",
            data_re_out => mul_re_out(593),
            data_im_out => mul_im_out(593)
        );

 
    UMUL_594 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(594),
            data_im_in => first_stage_im_out(594),
            re_multiplicator => "0011100001000010", --- 0.879028320312 + j-0.476806640625
            im_multiplicator => "1110000101111100",
            data_re_out => mul_re_out(594),
            data_im_out => mul_im_out(594)
        );

 
    UMUL_595 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(595),
            data_im_in => first_stage_im_out(595),
            re_multiplicator => "0011011101100101", --- 0.865539550781 + j-0.500915527344
            im_multiplicator => "1101111111110001",
            data_re_out => mul_re_out(595),
            data_im_out => mul_im_out(595)
        );

 
    UMUL_596 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(596),
            data_im_in => first_stage_im_out(596),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(596),
            data_im_out => mul_im_out(596)
        );

 
    UMUL_597 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(597),
            data_im_in => first_stage_im_out(597),
            re_multiplicator => "0011010110001010", --- 0.836547851562 + j-0.547912597656
            im_multiplicator => "1101110011101111",
            data_re_out => mul_re_out(597),
            data_im_out => mul_im_out(597)
        );

 
    UMUL_598 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(598),
            data_im_in => first_stage_im_out(598),
            re_multiplicator => "0011010010001101", --- 0.821105957031 + j-0.57080078125
            im_multiplicator => "1101101101111000",
            data_re_out => mul_re_out(598),
            data_im_out => mul_im_out(598)
        );

 
    UMUL_599 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(599),
            data_im_in => first_stage_im_out(599),
            re_multiplicator => "0011001110000110", --- 0.805053710938 + j-0.59326171875
            im_multiplicator => "1101101000001000",
            data_re_out => mul_re_out(599),
            data_im_out => mul_im_out(599)
        );

 
    UMUL_600 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(600),
            data_im_in => first_stage_im_out(600),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(600),
            data_im_out => mul_im_out(600)
        );

 
    UMUL_601 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(601),
            data_im_in => first_stage_im_out(601),
            re_multiplicator => "0011000101011001", --- 0.771057128906 + j-0.636779785156
            im_multiplicator => "1101011100111111",
            data_re_out => mul_re_out(601),
            data_im_out => mul_im_out(601)
        );

 
    UMUL_602 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(602),
            data_im_in => first_stage_im_out(602),
            re_multiplicator => "0011000000110100", --- 0.753173828125 + j-0.657836914062
            im_multiplicator => "1101010111100110",
            data_re_out => mul_re_out(602),
            data_im_out => mul_im_out(602)
        );

 
    UMUL_603 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(603),
            data_im_in => first_stage_im_out(603),
            re_multiplicator => "0010111100000110", --- 0.734741210938 + j-0.678344726562
            im_multiplicator => "1101010010010110",
            data_re_out => mul_re_out(603),
            data_im_out => mul_im_out(603)
        );

 
    UMUL_604 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(604),
            data_im_in => first_stage_im_out(604),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(604),
            data_im_out => mul_im_out(604)
        );

 
    UMUL_605 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(605),
            data_im_in => first_stage_im_out(605),
            re_multiplicator => "0010110010001110", --- 0.696166992188 + j-0.717895507812
            im_multiplicator => "1101001000001110",
            data_re_out => mul_re_out(605),
            data_im_out => mul_im_out(605)
        );

 
    UMUL_606 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(606),
            data_im_in => first_stage_im_out(606),
            re_multiplicator => "0010101101000101", --- 0.676086425781 + j-0.73681640625
            im_multiplicator => "1101000011011000",
            data_re_out => mul_re_out(606),
            data_im_out => mul_im_out(606)
        );

 
    UMUL_607 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(607),
            data_im_in => first_stage_im_out(607),
            re_multiplicator => "0010100111110100", --- 0.655517578125 + j-0.755187988281
            im_multiplicator => "1100111110101011",
            data_re_out => mul_re_out(607),
            data_im_out => mul_im_out(607)
        );

 
    UMUL_608 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(608),
            data_im_in => first_stage_im_out(608),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(608),
            data_im_out => mul_im_out(608)
        );

 
    UMUL_609 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(609),
            data_im_in => first_stage_im_out(609),
            re_multiplicator => "0010011100111000", --- 0.61279296875 + j-0.790222167969
            im_multiplicator => "1100110101101101",
            data_re_out => mul_re_out(609),
            data_im_out => mul_im_out(609)
        );

 
    UMUL_610 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(610),
            data_im_in => first_stage_im_out(610),
            re_multiplicator => "0010010111001111", --- 0.590759277344 + j-0.806823730469
            im_multiplicator => "1100110001011101",
            data_re_out => mul_re_out(610),
            data_im_out => mul_im_out(610)
        );

 
    UMUL_611 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(611),
            data_im_in => first_stage_im_out(611),
            re_multiplicator => "0010010001011110", --- 0.568237304688 + j-0.822875976562
            im_multiplicator => "1100101101010110",
            data_re_out => mul_re_out(611),
            data_im_out => mul_im_out(611)
        );

 
    UMUL_612 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(612),
            data_im_in => first_stage_im_out(612),
            re_multiplicator => "0010001011100111", --- 0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(612),
            data_im_out => mul_im_out(612)
        );

 
    UMUL_613 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(613),
            data_im_in => first_stage_im_out(613),
            re_multiplicator => "0010000101101000", --- 0.52197265625 + j-0.852966308594
            im_multiplicator => "1100100101101001",
            data_re_out => mul_re_out(613),
            data_im_out => mul_im_out(613)
        );

 
    UMUL_614 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(614),
            data_im_in => first_stage_im_out(614),
            re_multiplicator => "0001111111100011", --- 0.498229980469 + j-0.867065429688
            im_multiplicator => "1100100010000010",
            data_re_out => mul_re_out(614),
            data_im_out => mul_im_out(614)
        );

 
    UMUL_615 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(615),
            data_im_in => first_stage_im_out(615),
            re_multiplicator => "0001111001011000", --- 0.47412109375 + j-0.880493164062
            im_multiplicator => "1100011110100110",
            data_re_out => mul_re_out(615),
            data_im_out => mul_im_out(615)
        );

 
    UMUL_616 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(616),
            data_im_in => first_stage_im_out(616),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(616),
            data_im_out => mul_im_out(616)
        );

 
    UMUL_617 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(617),
            data_im_in => first_stage_im_out(617),
            re_multiplicator => "0001101100110000", --- 0.4248046875 + j-0.9052734375
            im_multiplicator => "1100011000010000",
            data_re_out => mul_re_out(617),
            data_im_out => mul_im_out(617)
        );

 
    UMUL_618 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(618),
            data_im_in => first_stage_im_out(618),
            re_multiplicator => "0001100110010011", --- 0.399597167969 + j-0.916687011719
            im_multiplicator => "1100010101010101",
            data_re_out => mul_re_out(618),
            data_im_out => mul_im_out(618)
        );

 
    UMUL_619 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(619),
            data_im_in => first_stage_im_out(619),
            re_multiplicator => "0001011111110010", --- 0.374145507812 + j-0.927368164062
            im_multiplicator => "1100010010100110",
            data_re_out => mul_re_out(619),
            data_im_out => mul_im_out(619)
        );

 
    UMUL_620 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(620),
            data_im_in => first_stage_im_out(620),
            re_multiplicator => "0001011001001100", --- 0.348388671875 + j-0.937316894531
            im_multiplicator => "1100010000000011",
            data_re_out => mul_re_out(620),
            data_im_out => mul_im_out(620)
        );

 
    UMUL_621 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(621),
            data_im_in => first_stage_im_out(621),
            re_multiplicator => "0001010010100010", --- 0.322387695312 + j-0.946594238281
            im_multiplicator => "1100001101101011",
            data_re_out => mul_re_out(621),
            data_im_out => mul_im_out(621)
        );

 
    UMUL_622 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(622),
            data_im_in => first_stage_im_out(622),
            re_multiplicator => "0001001011110100", --- 0.296142578125 + j-0.955139160156
            im_multiplicator => "1100001011011111",
            data_re_out => mul_re_out(622),
            data_im_out => mul_im_out(622)
        );

 
    UMUL_623 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(623),
            data_im_in => first_stage_im_out(623),
            re_multiplicator => "0001000101000010", --- 0.269653320312 + j-0.962951660156
            im_multiplicator => "1100001001011111",
            data_re_out => mul_re_out(623),
            data_im_out => mul_im_out(623)
        );

 
    UMUL_624 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(624),
            data_im_in => first_stage_im_out(624),
            re_multiplicator => "0000111110001101", --- 0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(624),
            data_im_out => mul_im_out(624)
        );

 
    UMUL_625 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(625),
            data_im_in => first_stage_im_out(625),
            re_multiplicator => "0000110111010101", --- 0.216125488281 + j-0.976379394531
            im_multiplicator => "1100000110000011",
            data_re_out => mul_re_out(625),
            data_im_out => mul_im_out(625)
        );

 
    UMUL_626 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(626),
            data_im_in => first_stage_im_out(626),
            re_multiplicator => "0000110000011010", --- 0.189086914062 + j-0.98193359375
            im_multiplicator => "1100000100101000",
            data_re_out => mul_re_out(626),
            data_im_out => mul_im_out(626)
        );

 
    UMUL_627 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(627),
            data_im_in => first_stage_im_out(627),
            re_multiplicator => "0000101001011100", --- 0.161865234375 + j-0.98681640625
            im_multiplicator => "1100000011011000",
            data_re_out => mul_re_out(627),
            data_im_out => mul_im_out(627)
        );

 
    UMUL_628 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(628),
            data_im_in => first_stage_im_out(628),
            re_multiplicator => "0000100010011101", --- 0.134582519531 + j-0.990905761719
            im_multiplicator => "1100000010010101",
            data_re_out => mul_re_out(628),
            data_im_out => mul_im_out(628)
        );

 
    UMUL_629 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(629),
            data_im_in => first_stage_im_out(629),
            re_multiplicator => "0000011011011100", --- 0.107177734375 + j-0.994262695312
            im_multiplicator => "1100000001011110",
            data_re_out => mul_re_out(629),
            data_im_out => mul_im_out(629)
        );

 
    UMUL_630 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(630),
            data_im_in => first_stage_im_out(630),
            re_multiplicator => "0000010100011010", --- 0.0797119140625 + j-0.996826171875
            im_multiplicator => "1100000000110100",
            data_re_out => mul_re_out(630),
            data_im_out => mul_im_out(630)
        );

 
    UMUL_631 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(631),
            data_im_in => first_stage_im_out(631),
            re_multiplicator => "0000001101010110", --- 0.0521240234375 + j-0.998657226562
            im_multiplicator => "1100000000010110",
            data_re_out => mul_re_out(631),
            data_im_out => mul_im_out(631)
        );

 
    UMUL_632 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(632),
            data_im_in => first_stage_im_out(632),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(632),
            data_im_out => mul_im_out(632)
        );

 
    UMUL_633 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(633),
            data_im_in => first_stage_im_out(633),
            re_multiplicator => "1111111111001110", --- -0.0030517578125 + j-1.0
            im_multiplicator => "1100000000000000",
            data_re_out => mul_re_out(633),
            data_im_out => mul_im_out(633)
        );

 
    UMUL_634 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(634),
            data_im_in => first_stage_im_out(634),
            re_multiplicator => "1111111000001001", --- -0.0307006835938 + j-0.99951171875
            im_multiplicator => "1100000000001000",
            data_re_out => mul_re_out(634),
            data_im_out => mul_im_out(634)
        );

 
    UMUL_635 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(635),
            data_im_in => first_stage_im_out(635),
            re_multiplicator => "1111110001000101", --- -0.0582885742188 + j-0.998291015625
            im_multiplicator => "1100000000011100",
            data_re_out => mul_re_out(635),
            data_im_out => mul_im_out(635)
        );

 
    UMUL_636 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(636),
            data_im_in => first_stage_im_out(636),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(636),
            data_im_out => mul_im_out(636)
        );

 
    UMUL_637 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(637),
            data_im_in => first_stage_im_out(637),
            re_multiplicator => "1111100011000000", --- -0.11328125 + j-0.993591308594
            im_multiplicator => "1100000001101001",
            data_re_out => mul_re_out(637),
            data_im_out => mul_im_out(637)
        );

 
    UMUL_638 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(638),
            data_im_in => first_stage_im_out(638),
            re_multiplicator => "1111011011111111", --- -0.140686035156 + j-0.990051269531
            im_multiplicator => "1100000010100011",
            data_re_out => mul_re_out(638),
            data_im_out => mul_im_out(638)
        );

 
    UMUL_639 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(639),
            data_im_in => first_stage_im_out(639),
            re_multiplicator => "1111010101000000", --- -0.16796875 + j-0.985778808594
            im_multiplicator => "1100000011101001",
            data_re_out => mul_re_out(639),
            data_im_out => mul_im_out(639)
        );

 
    UMUL_640 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(640),
            data_im_in => first_stage_im_out(640),
            data_re_out => mul_re_out(640),
            data_im_out => mul_im_out(640)
        );

 
    UMUL_641 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(641),
            data_im_in => first_stage_im_out(641),
            re_multiplicator => "0011111111111000", --- 0.99951171875 + j-0.0307006835938
            im_multiplicator => "1111111000001001",
            data_re_out => mul_re_out(641),
            data_im_out => mul_im_out(641)
        );

 
    UMUL_642 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(642),
            data_im_in => first_stage_im_out(642),
            re_multiplicator => "0011111111100001", --- 0.998107910156 + j-0.0613403320312
            im_multiplicator => "1111110000010011",
            data_re_out => mul_re_out(642),
            data_im_out => mul_im_out(642)
        );

 
    UMUL_643 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(643),
            data_im_in => first_stage_im_out(643),
            re_multiplicator => "0011111110111011", --- 0.995788574219 + j-0.0919189453125
            im_multiplicator => "1111101000011110",
            data_re_out => mul_re_out(643),
            data_im_out => mul_im_out(643)
        );

 
    UMUL_644 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(644),
            data_im_in => first_stage_im_out(644),
            re_multiplicator => "0011111110000101", --- 0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(644),
            data_im_out => mul_im_out(644)
        );

 
    UMUL_645 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(645),
            data_im_in => first_stage_im_out(645),
            re_multiplicator => "0011111101000000", --- 0.98828125 + j-0.152770996094
            im_multiplicator => "1111011000111001",
            data_re_out => mul_re_out(645),
            data_im_out => mul_im_out(645)
        );

 
    UMUL_646 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(646),
            data_im_in => first_stage_im_out(646),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(646),
            data_im_out => mul_im_out(646)
        );

 
    UMUL_647 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(647),
            data_im_in => first_stage_im_out(647),
            re_multiplicator => "0011111010001000", --- 0.97705078125 + j-0.213134765625
            im_multiplicator => "1111001001011100",
            data_re_out => mul_re_out(647),
            data_im_out => mul_im_out(647)
        );

 
    UMUL_648 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(648),
            data_im_in => first_stage_im_out(648),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(648),
            data_im_out => mul_im_out(648)
        );

 
    UMUL_649 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(649),
            data_im_in => first_stage_im_out(649),
            re_multiplicator => "0011110110010011", --- 0.962097167969 + j-0.272644042969
            im_multiplicator => "1110111010001101",
            data_re_out => mul_re_out(649),
            data_im_out => mul_im_out(649)
        );

 
    UMUL_650 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(650),
            data_im_in => first_stage_im_out(650),
            re_multiplicator => "0011110100000011", --- 0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(650),
            data_im_out => mul_im_out(650)
        );

 
    UMUL_651 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(651),
            data_im_in => first_stage_im_out(651),
            re_multiplicator => "0011110001100100", --- 0.943603515625 + j-0.331115722656
            im_multiplicator => "1110101011001111",
            data_re_out => mul_re_out(651),
            data_im_out => mul_im_out(651)
        );

 
    UMUL_652 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(652),
            data_im_in => first_stage_im_out(652),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(652),
            data_im_out => mul_im_out(652)
        );

 
    UMUL_653 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(653),
            data_im_in => first_stage_im_out(653),
            re_multiplicator => "0011101011111010", --- 0.921508789062 + j-0.388366699219
            im_multiplicator => "1110011100100101",
            data_re_out => mul_re_out(653),
            data_im_out => mul_im_out(653)
        );

 
    UMUL_654 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(654),
            data_im_in => first_stage_im_out(654),
            re_multiplicator => "0011101000110000", --- 0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(654),
            data_im_out => mul_im_out(654)
        );

 
    UMUL_655 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(655),
            data_im_in => first_stage_im_out(655),
            re_multiplicator => "0011100101011000", --- 0.89599609375 + j-0.444091796875
            im_multiplicator => "1110001110010100",
            data_re_out => mul_re_out(655),
            data_im_out => mul_im_out(655)
        );

 
    UMUL_656 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(656),
            data_im_in => first_stage_im_out(656),
            re_multiplicator => "0011100001110001", --- 0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(656),
            data_im_out => mul_im_out(656)
        );

 
    UMUL_657 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(657),
            data_im_in => first_stage_im_out(657),
            re_multiplicator => "0011011101111110", --- 0.867065429688 + j-0.498229980469
            im_multiplicator => "1110000000011101",
            data_re_out => mul_re_out(657),
            data_im_out => mul_im_out(657)
        );

 
    UMUL_658 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(658),
            data_im_in => first_stage_im_out(658),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(658),
            data_im_out => mul_im_out(658)
        );

 
    UMUL_659 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(659),
            data_im_in => first_stage_im_out(659),
            re_multiplicator => "0011010101101110", --- 0.834838867188 + j-0.550476074219
            im_multiplicator => "1101110011000101",
            data_re_out => mul_re_out(659),
            data_im_out => mul_im_out(659)
        );

 
    UMUL_660 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(660),
            data_im_in => first_stage_im_out(660),
            re_multiplicator => "0011010001010011", --- 0.817565917969 + j-0.575805664062
            im_multiplicator => "1101101100100110",
            data_re_out => mul_re_out(660),
            data_im_out => mul_im_out(660)
        );

 
    UMUL_661 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(661),
            data_im_in => first_stage_im_out(661),
            re_multiplicator => "0011001100101100", --- 0.799560546875 + j-0.600646972656
            im_multiplicator => "1101100110001111",
            data_re_out => mul_re_out(661),
            data_im_out => mul_im_out(661)
        );

 
    UMUL_662 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(662),
            data_im_in => first_stage_im_out(662),
            re_multiplicator => "0011000111111000", --- 0.78076171875 + j-0.624877929688
            im_multiplicator => "1101100000000010",
            data_re_out => mul_re_out(662),
            data_im_out => mul_im_out(662)
        );

 
    UMUL_663 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(663),
            data_im_in => first_stage_im_out(663),
            re_multiplicator => "0011000010111000", --- 0.76123046875 + j-0.648498535156
            im_multiplicator => "1101011001111111",
            data_re_out => mul_re_out(663),
            data_im_out => mul_im_out(663)
        );

 
    UMUL_664 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(664),
            data_im_in => first_stage_im_out(664),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(664),
            data_im_out => mul_im_out(664)
        );

 
    UMUL_665 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(665),
            data_im_in => first_stage_im_out(665),
            re_multiplicator => "0010111000010101", --- 0.720031738281 + j-0.693969726562
            im_multiplicator => "1101001110010110",
            data_re_out => mul_re_out(665),
            data_im_out => mul_im_out(665)
        );

 
    UMUL_666 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(666),
            data_im_in => first_stage_im_out(666),
            re_multiplicator => "0010110010110010", --- 0.698364257812 + j-0.715759277344
            im_multiplicator => "1101001000110001",
            data_re_out => mul_re_out(666),
            data_im_out => mul_im_out(666)
        );

 
    UMUL_667 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(667),
            data_im_in => first_stage_im_out(667),
            re_multiplicator => "0010101101000101", --- 0.676086425781 + j-0.73681640625
            im_multiplicator => "1101000011011000",
            data_re_out => mul_re_out(667),
            data_im_out => mul_im_out(667)
        );

 
    UMUL_668 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(668),
            data_im_in => first_stage_im_out(668),
            re_multiplicator => "0010100111001110", --- 0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(668),
            data_im_out => mul_im_out(668)
        );

 
    UMUL_669 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(669),
            data_im_in => first_stage_im_out(669),
            re_multiplicator => "0010100001001100", --- 0.629638671875 + j-0.776916503906
            im_multiplicator => "1100111001000111",
            data_re_out => mul_re_out(669),
            data_im_out => mul_im_out(669)
        );

 
    UMUL_670 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(670),
            data_im_in => first_stage_im_out(670),
            re_multiplicator => "0010011011000001", --- 0.605529785156 + j-0.795837402344
            im_multiplicator => "1100110100010001",
            data_re_out => mul_re_out(670),
            data_im_out => mul_im_out(670)
        );

 
    UMUL_671 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(671),
            data_im_in => first_stage_im_out(671),
            re_multiplicator => "0010010100101100", --- 0.580810546875 + j-0.814025878906
            im_multiplicator => "1100101111100111",
            data_re_out => mul_re_out(671),
            data_im_out => mul_im_out(671)
        );

 
    UMUL_672 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(672),
            data_im_in => first_stage_im_out(672),
            re_multiplicator => "0010001110001110", --- 0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(672),
            data_im_out => mul_im_out(672)
        );

 
    UMUL_673 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(673),
            data_im_in => first_stage_im_out(673),
            re_multiplicator => "0010000111101000", --- 0.52978515625 + j-0.84814453125
            im_multiplicator => "1100100110111000",
            data_re_out => mul_re_out(673),
            data_im_out => mul_im_out(673)
        );

 
    UMUL_674 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(674),
            data_im_in => first_stage_im_out(674),
            re_multiplicator => "0010000000111010", --- 0.503540039062 + j-0.863952636719
            im_multiplicator => "1100100010110101",
            data_re_out => mul_re_out(674),
            data_im_out => mul_im_out(674)
        );

 
    UMUL_675 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(675),
            data_im_in => first_stage_im_out(675),
            re_multiplicator => "0001111010000100", --- 0.476806640625 + j-0.879028320312
            im_multiplicator => "1100011110111110",
            data_re_out => mul_re_out(675),
            data_im_out => mul_im_out(675)
        );

 
    UMUL_676 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(676),
            data_im_in => first_stage_im_out(676),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(676),
            data_im_out => mul_im_out(676)
        );

 
    UMUL_677 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(677),
            data_im_in => first_stage_im_out(677),
            re_multiplicator => "0001101100000010", --- 0.421997070312 + j-0.906616210938
            im_multiplicator => "1100010111111010",
            data_re_out => mul_re_out(677),
            data_im_out => mul_im_out(677)
        );

 
    UMUL_678 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(678),
            data_im_in => first_stage_im_out(678),
            re_multiplicator => "0001100100110111", --- 0.393981933594 + j-0.919128417969
            im_multiplicator => "1100010100101101",
            data_re_out => mul_re_out(678),
            data_im_out => mul_im_out(678)
        );

 
    UMUL_679 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(679),
            data_im_in => first_stage_im_out(679),
            re_multiplicator => "0001011101100110", --- 0.365600585938 + j-0.930786132812
            im_multiplicator => "1100010001101110",
            data_re_out => mul_re_out(679),
            data_im_out => mul_im_out(679)
        );

 
    UMUL_680 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(680),
            data_im_in => first_stage_im_out(680),
            re_multiplicator => "0001010110010000", --- 0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(680),
            data_im_out => mul_im_out(680)
        );

 
    UMUL_681 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(681),
            data_im_in => first_stage_im_out(681),
            re_multiplicator => "0001001110110100", --- 0.307861328125 + j-0.951416015625
            im_multiplicator => "1100001100011100",
            data_re_out => mul_re_out(681),
            data_im_out => mul_im_out(681)
        );

 
    UMUL_682 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(682),
            data_im_in => first_stage_im_out(682),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(682),
            data_im_out => mul_im_out(682)
        );

 
    UMUL_683 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(683),
            data_im_in => first_stage_im_out(683),
            re_multiplicator => "0000111111101110", --- 0.248901367188 + j-0.968505859375
            im_multiplicator => "1100001000000100",
            data_re_out => mul_re_out(683),
            data_im_out => mul_im_out(683)
        );

 
    UMUL_684 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(684),
            data_im_in => first_stage_im_out(684),
            re_multiplicator => "0000111000000110", --- 0.219116210938 + j-0.975708007812
            im_multiplicator => "1100000110001110",
            data_re_out => mul_re_out(684),
            data_im_out => mul_im_out(684)
        );

 
    UMUL_685 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(685),
            data_im_in => first_stage_im_out(685),
            re_multiplicator => "0000110000011010", --- 0.189086914062 + j-0.98193359375
            im_multiplicator => "1100000100101000",
            data_re_out => mul_re_out(685),
            data_im_out => mul_im_out(685)
        );

 
    UMUL_686 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(686),
            data_im_in => first_stage_im_out(686),
            re_multiplicator => "0000101000101011", --- 0.158874511719 + j-0.9873046875
            im_multiplicator => "1100000011010000",
            data_re_out => mul_re_out(686),
            data_im_out => mul_im_out(686)
        );

 
    UMUL_687 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(687),
            data_im_in => first_stage_im_out(687),
            re_multiplicator => "0000100000111001", --- 0.128479003906 + j-0.99169921875
            im_multiplicator => "1100000010001000",
            data_re_out => mul_re_out(687),
            data_im_out => mul_im_out(687)
        );

 
    UMUL_688 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(688),
            data_im_in => first_stage_im_out(688),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(688),
            data_im_out => mul_im_out(688)
        );

 
    UMUL_689 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(689),
            data_im_in => first_stage_im_out(689),
            re_multiplicator => "0000010001010001", --- 0.0674438476562 + j-0.997741699219
            im_multiplicator => "1100000000100101",
            data_re_out => mul_re_out(689),
            data_im_out => mul_im_out(689)
        );

 
    UMUL_690 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(690),
            data_im_in => first_stage_im_out(690),
            re_multiplicator => "0000001001011011", --- 0.0368041992188 + j-0.999328613281
            im_multiplicator => "1100000000001011",
            data_re_out => mul_re_out(690),
            data_im_out => mul_im_out(690)
        );

 
    UMUL_691 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(691),
            data_im_in => first_stage_im_out(691),
            re_multiplicator => "0000000001100101", --- 0.00616455078125 + j-1.0
            im_multiplicator => "1100000000000000",
            data_re_out => mul_re_out(691),
            data_im_out => mul_im_out(691)
        );

 
    UMUL_692 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(692),
            data_im_in => first_stage_im_out(692),
            re_multiplicator => "1111111001101110", --- -0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(692),
            data_im_out => mul_im_out(692)
        );

 
    UMUL_693 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(693),
            data_im_in => first_stage_im_out(693),
            re_multiplicator => "1111110001111000", --- -0.05517578125 + j-0.998474121094
            im_multiplicator => "1100000000011001",
            data_re_out => mul_re_out(693),
            data_im_out => mul_im_out(693)
        );

 
    UMUL_694 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(694),
            data_im_in => first_stage_im_out(694),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(694),
            data_im_out => mul_im_out(694)
        );

 
    UMUL_695 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(695),
            data_im_in => first_stage_im_out(695),
            re_multiplicator => "1111100010001110", --- -0.116333007812 + j-0.993225097656
            im_multiplicator => "1100000001101111",
            data_re_out => mul_re_out(695),
            data_im_out => mul_im_out(695)
        );

 
    UMUL_696 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(696),
            data_im_in => first_stage_im_out(696),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(696),
            data_im_out => mul_im_out(696)
        );

 
    UMUL_697 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(697),
            data_im_in => first_stage_im_out(697),
            re_multiplicator => "1111010010101100", --- -0.177001953125 + j-0.984191894531
            im_multiplicator => "1100000100000011",
            data_re_out => mul_re_out(697),
            data_im_out => mul_im_out(697)
        );

 
    UMUL_698 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(698),
            data_im_in => first_stage_im_out(698),
            re_multiplicator => "1111001010111111", --- -0.207092285156 + j-0.978332519531
            im_multiplicator => "1100000101100011",
            data_re_out => mul_re_out(698),
            data_im_out => mul_im_out(698)
        );

 
    UMUL_699 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(699),
            data_im_in => first_stage_im_out(699),
            re_multiplicator => "1111000011010101", --- -0.236999511719 + j-0.971496582031
            im_multiplicator => "1100000111010011",
            data_re_out => mul_re_out(699),
            data_im_out => mul_im_out(699)
        );

 
    UMUL_700 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(700),
            data_im_in => first_stage_im_out(700),
            re_multiplicator => "1110111011101110", --- -0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(700),
            data_im_out => mul_im_out(700)
        );

 
    UMUL_701 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(701),
            data_im_in => first_stage_im_out(701),
            re_multiplicator => "1110110100001100", --- -0.296142578125 + j-0.955139160156
            im_multiplicator => "1100001011011111",
            data_re_out => mul_re_out(701),
            data_im_out => mul_im_out(701)
        );

 
    UMUL_702 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(702),
            data_im_in => first_stage_im_out(702),
            re_multiplicator => "1110101100101110", --- -0.325317382812 + j-0.945617675781
            im_multiplicator => "1100001101111011",
            data_re_out => mul_re_out(702),
            data_im_out => mul_im_out(702)
        );

 
    UMUL_703 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(703),
            data_im_in => first_stage_im_out(703),
            re_multiplicator => "1110100101010101", --- -0.354187011719 + j-0.935180664062
            im_multiplicator => "1100010000100110",
            data_re_out => mul_re_out(703),
            data_im_out => mul_im_out(703)
        );

 
    UMUL_704 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(704),
            data_im_in => first_stage_im_out(704),
            data_re_out => mul_re_out(704),
            data_im_out => mul_im_out(704)
        );

 
    UMUL_705 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(705),
            data_im_in => first_stage_im_out(705),
            re_multiplicator => "0011111111110111", --- 0.999450683594 + j-0.0337524414062
            im_multiplicator => "1111110111010111",
            data_re_out => mul_re_out(705),
            data_im_out => mul_im_out(705)
        );

 
    UMUL_706 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(706),
            data_im_in => first_stage_im_out(706),
            re_multiplicator => "0011111111011011", --- 0.997741699219 + j-0.0674438476562
            im_multiplicator => "1111101110101111",
            data_re_out => mul_re_out(706),
            data_im_out => mul_im_out(706)
        );

 
    UMUL_707 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(707),
            data_im_in => first_stage_im_out(707),
            re_multiplicator => "0011111110101100", --- 0.994873046875 + j-0.10107421875
            im_multiplicator => "1111100110001000",
            data_re_out => mul_re_out(707),
            data_im_out => mul_im_out(707)
        );

 
    UMUL_708 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(708),
            data_im_in => first_stage_im_out(708),
            re_multiplicator => "0011111101101011", --- 0.990905761719 + j-0.134582519531
            im_multiplicator => "1111011101100011",
            data_re_out => mul_re_out(708),
            data_im_out => mul_im_out(708)
        );

 
    UMUL_709 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(709),
            data_im_in => first_stage_im_out(709),
            re_multiplicator => "0011111100010111", --- 0.985778808594 + j-0.16796875
            im_multiplicator => "1111010101000000",
            data_re_out => mul_re_out(709),
            data_im_out => mul_im_out(709)
        );

 
    UMUL_710 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(710),
            data_im_in => first_stage_im_out(710),
            re_multiplicator => "0011111010110001", --- 0.979553222656 + j-0.201110839844
            im_multiplicator => "1111001100100001",
            data_re_out => mul_re_out(710),
            data_im_out => mul_im_out(710)
        );

 
    UMUL_711 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(711),
            data_im_in => first_stage_im_out(711),
            re_multiplicator => "0011111000111001", --- 0.972229003906 + j-0.234069824219
            im_multiplicator => "1111000100000101",
            data_re_out => mul_re_out(711),
            data_im_out => mul_im_out(711)
        );

 
    UMUL_712 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(712),
            data_im_in => first_stage_im_out(712),
            re_multiplicator => "0011110110101111", --- 0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(712),
            data_im_out => mul_im_out(712)
        );

 
    UMUL_713 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(713),
            data_im_in => first_stage_im_out(713),
            re_multiplicator => "0011110100010010", --- 0.954223632812 + j-0.299072265625
            im_multiplicator => "1110110011011100",
            data_re_out => mul_re_out(713),
            data_im_out => mul_im_out(713)
        );

 
    UMUL_714 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(714),
            data_im_in => first_stage_im_out(714),
            re_multiplicator => "0011110001100100", --- 0.943603515625 + j-0.331115722656
            im_multiplicator => "1110101011001111",
            data_re_out => mul_re_out(714),
            data_im_out => mul_im_out(714)
        );

 
    UMUL_715 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(715),
            data_im_in => first_stage_im_out(715),
            re_multiplicator => "0011101110100100", --- 0.931884765625 + j-0.362731933594
            im_multiplicator => "1110100011001001",
            data_re_out => mul_re_out(715),
            data_im_out => mul_im_out(715)
        );

 
    UMUL_716 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(716),
            data_im_in => first_stage_im_out(716),
            re_multiplicator => "0011101011010011", --- 0.919128417969 + j-0.393981933594
            im_multiplicator => "1110011011001001",
            data_re_out => mul_re_out(716),
            data_im_out => mul_im_out(716)
        );

 
    UMUL_717 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(717),
            data_im_in => first_stage_im_out(717),
            re_multiplicator => "0011100111110000", --- 0.9052734375 + j-0.4248046875
            im_multiplicator => "1110010011010000",
            data_re_out => mul_re_out(717),
            data_im_out => mul_im_out(717)
        );

 
    UMUL_718 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(718),
            data_im_in => first_stage_im_out(718),
            re_multiplicator => "0011100011111101", --- 0.890441894531 + j-0.455078125
            im_multiplicator => "1110001011100000",
            data_re_out => mul_re_out(718),
            data_im_out => mul_im_out(718)
        );

 
    UMUL_719 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(719),
            data_im_in => first_stage_im_out(719),
            re_multiplicator => "0011011111111001", --- 0.874572753906 + j-0.48486328125
            im_multiplicator => "1110000011111000",
            data_re_out => mul_re_out(719),
            data_im_out => mul_im_out(719)
        );

 
    UMUL_720 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(720),
            data_im_in => first_stage_im_out(720),
            re_multiplicator => "0011011011100101", --- 0.857727050781 + j-0.514099121094
            im_multiplicator => "1101111100011001",
            data_re_out => mul_re_out(720),
            data_im_out => mul_im_out(720)
        );

 
    UMUL_721 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(721),
            data_im_in => first_stage_im_out(721),
            re_multiplicator => "0011010111000001", --- 0.839904785156 + j-0.542724609375
            im_multiplicator => "1101110101000100",
            data_re_out => mul_re_out(721),
            data_im_out => mul_im_out(721)
        );

 
    UMUL_722 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(722),
            data_im_in => first_stage_im_out(722),
            re_multiplicator => "0011010010001101", --- 0.821105957031 + j-0.57080078125
            im_multiplicator => "1101101101111000",
            data_re_out => mul_re_out(722),
            data_im_out => mul_im_out(722)
        );

 
    UMUL_723 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(723),
            data_im_in => first_stage_im_out(723),
            re_multiplicator => "0011001101001010", --- 0.801391601562 + j-0.59814453125
            im_multiplicator => "1101100110111000",
            data_re_out => mul_re_out(723),
            data_im_out => mul_im_out(723)
        );

 
    UMUL_724 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(724),
            data_im_in => first_stage_im_out(724),
            re_multiplicator => "0011000111111000", --- 0.78076171875 + j-0.624877929688
            im_multiplicator => "1101100000000010",
            data_re_out => mul_re_out(724),
            data_im_out => mul_im_out(724)
        );

 
    UMUL_725 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(725),
            data_im_in => first_stage_im_out(725),
            re_multiplicator => "0011000010010111", --- 0.759216308594 + j-0.650817871094
            im_multiplicator => "1101011001011001",
            data_re_out => mul_re_out(725),
            data_im_out => mul_im_out(725)
        );

 
    UMUL_726 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(726),
            data_im_in => first_stage_im_out(726),
            re_multiplicator => "0010111100101000", --- 0.73681640625 + j-0.676086425781
            im_multiplicator => "1101010010111011",
            data_re_out => mul_re_out(726),
            data_im_out => mul_im_out(726)
        );

 
    UMUL_727 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(727),
            data_im_in => first_stage_im_out(727),
            re_multiplicator => "0010110110101011", --- 0.713562011719 + j-0.700561523438
            im_multiplicator => "1101001100101010",
            data_re_out => mul_re_out(727),
            data_im_out => mul_im_out(727)
        );

 
    UMUL_728 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(728),
            data_im_in => first_stage_im_out(728),
            re_multiplicator => "0010110000100001", --- 0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(728),
            data_im_out => mul_im_out(728)
        );

 
    UMUL_729 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(729),
            data_im_in => first_stage_im_out(729),
            re_multiplicator => "0010101010001011", --- 0.664733886719 + j-0.7470703125
            im_multiplicator => "1101000000110000",
            data_re_out => mul_re_out(729),
            data_im_out => mul_im_out(729)
        );

 
    UMUL_730 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(730),
            data_im_in => first_stage_im_out(730),
            re_multiplicator => "0010100011100111", --- 0.639099121094 + j-0.769104003906
            im_multiplicator => "1100111011000111",
            data_re_out => mul_re_out(730),
            data_im_out => mul_im_out(730)
        );

 
    UMUL_731 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(731),
            data_im_in => first_stage_im_out(731),
            re_multiplicator => "0010011100111000", --- 0.61279296875 + j-0.790222167969
            im_multiplicator => "1100110101101101",
            data_re_out => mul_re_out(731),
            data_im_out => mul_im_out(731)
        );

 
    UMUL_732 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(732),
            data_im_in => first_stage_im_out(732),
            re_multiplicator => "0010010101111110", --- 0.585815429688 + j-0.810485839844
            im_multiplicator => "1100110000100001",
            data_re_out => mul_re_out(732),
            data_im_out => mul_im_out(732)
        );

 
    UMUL_733 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(733),
            data_im_in => first_stage_im_out(733),
            re_multiplicator => "0010001110111000", --- 0.55810546875 + j-0.829772949219
            im_multiplicator => "1100101011100101",
            data_re_out => mul_re_out(733),
            data_im_out => mul_im_out(733)
        );

 
    UMUL_734 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(734),
            data_im_in => first_stage_im_out(734),
            re_multiplicator => "0010000111101000", --- 0.52978515625 + j-0.84814453125
            im_multiplicator => "1100100110111000",
            data_re_out => mul_re_out(734),
            data_im_out => mul_im_out(734)
        );

 
    UMUL_735 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(735),
            data_im_in => first_stage_im_out(735),
            re_multiplicator => "0010000000001111", --- 0.500915527344 + j-0.865539550781
            im_multiplicator => "1100100010011011",
            data_re_out => mul_re_out(735),
            data_im_out => mul_im_out(735)
        );

 
    UMUL_736 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(736),
            data_im_in => first_stage_im_out(736),
            re_multiplicator => "0001111000101011", --- 0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(736),
            data_im_out => mul_im_out(736)
        );

 
    UMUL_737 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(737),
            data_im_in => first_stage_im_out(737),
            re_multiplicator => "0001110000111111", --- 0.441345214844 + j-0.897338867188
            im_multiplicator => "1100011010010010",
            data_re_out => mul_re_out(737),
            data_im_out => mul_im_out(737)
        );

 
    UMUL_738 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(738),
            data_im_in => first_stage_im_out(738),
            re_multiplicator => "0001101001001011", --- 0.410827636719 + j-0.911682128906
            im_multiplicator => "1100010110100111",
            data_re_out => mul_re_out(738),
            data_im_out => mul_im_out(738)
        );

 
    UMUL_739 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(739),
            data_im_in => first_stage_im_out(739),
            re_multiplicator => "0001100001001111", --- 0.379821777344 + j-0.925048828125
            im_multiplicator => "1100010011001100",
            data_re_out => mul_re_out(739),
            data_im_out => mul_im_out(739)
        );

 
    UMUL_740 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(740),
            data_im_in => first_stage_im_out(740),
            re_multiplicator => "0001011001001100", --- 0.348388671875 + j-0.937316894531
            im_multiplicator => "1100010000000011",
            data_re_out => mul_re_out(740),
            data_im_out => mul_im_out(740)
        );

 
    UMUL_741 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(741),
            data_im_in => first_stage_im_out(741),
            re_multiplicator => "0001010001000011", --- 0.316589355469 + j-0.948547363281
            im_multiplicator => "1100001101001011",
            data_re_out => mul_re_out(741),
            data_im_out => mul_im_out(741)
        );

 
    UMUL_742 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(742),
            data_im_in => first_stage_im_out(742),
            re_multiplicator => "0001001000110100", --- 0.284423828125 + j-0.958679199219
            im_multiplicator => "1100001010100101",
            data_re_out => mul_re_out(742),
            data_im_out => mul_im_out(742)
        );

 
    UMUL_743 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(743),
            data_im_in => first_stage_im_out(743),
            re_multiplicator => "0001000000011111", --- 0.251892089844 + j-0.9677734375
            im_multiplicator => "1100001000010000",
            data_re_out => mul_re_out(743),
            data_im_out => mul_im_out(743)
        );

 
    UMUL_744 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(744),
            data_im_in => first_stage_im_out(744),
            re_multiplicator => "0000111000000110", --- 0.219116210938 + j-0.975708007812
            im_multiplicator => "1100000110001110",
            data_re_out => mul_re_out(744),
            data_im_out => mul_im_out(744)
        );

 
    UMUL_745 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(745),
            data_im_in => first_stage_im_out(745),
            re_multiplicator => "0000101111101000", --- 0.18603515625 + j-0.982543945312
            im_multiplicator => "1100000100011110",
            data_re_out => mul_re_out(745),
            data_im_out => mul_im_out(745)
        );

 
    UMUL_746 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(746),
            data_im_in => first_stage_im_out(746),
            re_multiplicator => "0000100111000111", --- 0.152770996094 + j-0.98828125
            im_multiplicator => "1100000011000000",
            data_re_out => mul_re_out(746),
            data_im_out => mul_im_out(746)
        );

 
    UMUL_747 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(747),
            data_im_in => first_stage_im_out(747),
            re_multiplicator => "0000011110100100", --- 0.119384765625 + j-0.992858886719
            im_multiplicator => "1100000001110101",
            data_re_out => mul_re_out(747),
            data_im_out => mul_im_out(747)
        );

 
    UMUL_748 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(748),
            data_im_in => first_stage_im_out(748),
            re_multiplicator => "0000010101111110", --- 0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(748),
            data_im_out => mul_im_out(748)
        );

 
    UMUL_749 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(749),
            data_im_in => first_stage_im_out(749),
            re_multiplicator => "0000001101010110", --- 0.0521240234375 + j-0.998657226562
            im_multiplicator => "1100000000010110",
            data_re_out => mul_re_out(749),
            data_im_out => mul_im_out(749)
        );

 
    UMUL_750 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(750),
            data_im_in => first_stage_im_out(750),
            re_multiplicator => "0000000100101110", --- 0.0184326171875 + j-0.999816894531
            im_multiplicator => "1100000000000011",
            data_re_out => mul_re_out(750),
            data_im_out => mul_im_out(750)
        );

 
    UMUL_751 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(751),
            data_im_in => first_stage_im_out(751),
            re_multiplicator => "1111111100000101", --- -0.0153198242188 + j-0.999877929688
            im_multiplicator => "1100000000000010",
            data_re_out => mul_re_out(751),
            data_im_out => mul_im_out(751)
        );

 
    UMUL_752 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(752),
            data_im_in => first_stage_im_out(752),
            re_multiplicator => "1111110011011100", --- -0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(752),
            data_im_out => mul_im_out(752)
        );

 
    UMUL_753 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(753),
            data_im_in => first_stage_im_out(753),
            re_multiplicator => "1111101010110100", --- -0.082763671875 + j-0.99658203125
            im_multiplicator => "1100000000111000",
            data_re_out => mul_re_out(753),
            data_im_out => mul_im_out(753)
        );

 
    UMUL_754 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(754),
            data_im_in => first_stage_im_out(754),
            re_multiplicator => "1111100010001110", --- -0.116333007812 + j-0.993225097656
            im_multiplicator => "1100000001101111",
            data_re_out => mul_re_out(754),
            data_im_out => mul_im_out(754)
        );

 
    UMUL_755 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(755),
            data_im_in => first_stage_im_out(755),
            re_multiplicator => "1111011001101010", --- -0.149780273438 + j-0.988708496094
            im_multiplicator => "1100000010111001",
            data_re_out => mul_re_out(755),
            data_im_out => mul_im_out(755)
        );

 
    UMUL_756 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(756),
            data_im_in => first_stage_im_out(756),
            re_multiplicator => "1111010001001001", --- -0.183044433594 + j-0.983093261719
            im_multiplicator => "1100000100010101",
            data_re_out => mul_re_out(756),
            data_im_out => mul_im_out(756)
        );

 
    UMUL_757 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(757),
            data_im_in => first_stage_im_out(757),
            re_multiplicator => "1111001000101011", --- -0.216125488281 + j-0.976379394531
            im_multiplicator => "1100000110000011",
            data_re_out => mul_re_out(757),
            data_im_out => mul_im_out(757)
        );

 
    UMUL_758 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(758),
            data_im_in => first_stage_im_out(758),
            re_multiplicator => "1111000000010010", --- -0.248901367188 + j-0.968505859375
            im_multiplicator => "1100001000000100",
            data_re_out => mul_re_out(758),
            data_im_out => mul_im_out(758)
        );

 
    UMUL_759 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(759),
            data_im_in => first_stage_im_out(759),
            re_multiplicator => "1110110111111100", --- -0.281494140625 + j-0.959594726562
            im_multiplicator => "1100001010010110",
            data_re_out => mul_re_out(759),
            data_im_out => mul_im_out(759)
        );

 
    UMUL_760 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(760),
            data_im_in => first_stage_im_out(760),
            re_multiplicator => "1110101111101101", --- -0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(760),
            data_im_out => mul_im_out(760)
        );

 
    UMUL_761 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(761),
            data_im_in => first_stage_im_out(761),
            re_multiplicator => "1110100111100011", --- -0.345520019531 + j-0.938415527344
            im_multiplicator => "1100001111110001",
            data_re_out => mul_re_out(761),
            data_im_out => mul_im_out(761)
        );

 
    UMUL_762 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(762),
            data_im_in => first_stage_im_out(762),
            re_multiplicator => "1110011111011111", --- -0.377014160156 + j-0.926208496094
            im_multiplicator => "1100010010111001",
            data_re_out => mul_re_out(762),
            data_im_out => mul_im_out(762)
        );

 
    UMUL_763 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(763),
            data_im_in => first_stage_im_out(763),
            re_multiplicator => "1110010111100011", --- -0.408020019531 + j-0.912963867188
            im_multiplicator => "1100010110010010",
            data_re_out => mul_re_out(763),
            data_im_out => mul_im_out(763)
        );

 
    UMUL_764 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(764),
            data_im_in => first_stage_im_out(764),
            re_multiplicator => "1110001111101110", --- -0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(764),
            data_im_out => mul_im_out(764)
        );

 
    UMUL_765 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(765),
            data_im_in => first_stage_im_out(765),
            re_multiplicator => "1110001000000001", --- -0.468688964844 + j-0.883361816406
            im_multiplicator => "1100011101110111",
            data_re_out => mul_re_out(765),
            data_im_out => mul_im_out(765)
        );

 
    UMUL_766 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(766),
            data_im_in => first_stage_im_out(766),
            re_multiplicator => "1110000000011101", --- -0.498229980469 + j-0.867065429688
            im_multiplicator => "1100100010000010",
            data_re_out => mul_re_out(766),
            data_im_out => mul_im_out(766)
        );

 
    UMUL_767 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(767),
            data_im_in => first_stage_im_out(767),
            re_multiplicator => "1101111001000010", --- -0.527221679688 + j-0.849731445312
            im_multiplicator => "1100100110011110",
            data_re_out => mul_re_out(767),
            data_im_out => mul_im_out(767)
        );

 
    UMUL_768 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(768),
            data_im_in => first_stage_im_out(768),
            data_re_out => mul_re_out(768),
            data_im_out => mul_im_out(768)
        );

 
    UMUL_769 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(769),
            data_im_in => first_stage_im_out(769),
            re_multiplicator => "0011111111110101", --- 0.999328613281 + j-0.0368041992188
            im_multiplicator => "1111110110100101",
            data_re_out => mul_re_out(769),
            data_im_out => mul_im_out(769)
        );

 
    UMUL_770 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(770),
            data_im_in => first_stage_im_out(770),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(770),
            data_im_out => mul_im_out(770)
        );

 
    UMUL_771 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(771),
            data_im_in => first_stage_im_out(771),
            re_multiplicator => "0011111110011100", --- 0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(771),
            data_im_out => mul_im_out(771)
        );

 
    UMUL_772 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(772),
            data_im_in => first_stage_im_out(772),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(772),
            data_im_out => mul_im_out(772)
        );

 
    UMUL_773 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(773),
            data_im_in => first_stage_im_out(773),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(773),
            data_im_out => mul_im_out(773)
        );

 
    UMUL_774 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(774),
            data_im_in => first_stage_im_out(774),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(774),
            data_im_out => mul_im_out(774)
        );

 
    UMUL_775 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(775),
            data_im_in => first_stage_im_out(775),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(775),
            data_im_out => mul_im_out(775)
        );

 
    UMUL_776 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(776),
            data_im_in => first_stage_im_out(776),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(776),
            data_im_out => mul_im_out(776)
        );

 
    UMUL_777 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(777),
            data_im_in => first_stage_im_out(777),
            re_multiplicator => "0011110010000101", --- 0.945617675781 + j-0.325317382812
            im_multiplicator => "1110101100101110",
            data_re_out => mul_re_out(777),
            data_im_out => mul_im_out(777)
        );

 
    UMUL_778 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(778),
            data_im_in => first_stage_im_out(778),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(778),
            data_im_out => mul_im_out(778)
        );

 
    UMUL_779 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(779),
            data_im_in => first_stage_im_out(779),
            re_multiplicator => "0011101011010011", --- 0.919128417969 + j-0.393981933594
            im_multiplicator => "1110011011001001",
            data_re_out => mul_re_out(779),
            data_im_out => mul_im_out(779)
        );

 
    UMUL_780 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(780),
            data_im_in => first_stage_im_out(780),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(780),
            data_im_out => mul_im_out(780)
        );

 
    UMUL_781 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(781),
            data_im_in => first_stage_im_out(781),
            re_multiplicator => "0011100011001111", --- 0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(781),
            data_im_out => mul_im_out(781)
        );

 
    UMUL_782 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(782),
            data_im_in => first_stage_im_out(782),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(782),
            data_im_out => mul_im_out(782)
        );

 
    UMUL_783 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(783),
            data_im_in => first_stage_im_out(783),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(783),
            data_im_out => mul_im_out(783)
        );

 
    UMUL_784 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(784),
            data_im_in => first_stage_im_out(784),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(784),
            data_im_out => mul_im_out(784)
        );

 
    UMUL_785 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(785),
            data_im_in => first_stage_im_out(785),
            re_multiplicator => "0011001111011111", --- 0.810485839844 + j-0.585815429688
            im_multiplicator => "1101101010000010",
            data_re_out => mul_re_out(785),
            data_im_out => mul_im_out(785)
        );

 
    UMUL_786 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(786),
            data_im_in => first_stage_im_out(786),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(786),
            data_im_out => mul_im_out(786)
        );

 
    UMUL_787 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(787),
            data_im_in => first_stage_im_out(787),
            re_multiplicator => "0011000011111001", --- 0.765197753906 + j-0.643859863281
            im_multiplicator => "1101011011001011",
            data_re_out => mul_re_out(787),
            data_im_out => mul_im_out(787)
        );

 
    UMUL_788 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(788),
            data_im_in => first_stage_im_out(788),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(788),
            data_im_out => mul_im_out(788)
        );

 
    UMUL_789 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(789),
            data_im_in => first_stage_im_out(789),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(789),
            data_im_out => mul_im_out(789)
        );

 
    UMUL_790 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(790),
            data_im_in => first_stage_im_out(790),
            re_multiplicator => "0010110000100001", --- 0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(790),
            data_im_out => mul_im_out(790)
        );

 
    UMUL_791 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(791),
            data_im_in => first_stage_im_out(791),
            re_multiplicator => "0010101001100101", --- 0.662414550781 + j-0.749145507812
            im_multiplicator => "1101000000001110",
            data_re_out => mul_re_out(791),
            data_im_out => mul_im_out(791)
        );

 
    UMUL_792 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(792),
            data_im_in => first_stage_im_out(792),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(792),
            data_im_out => mul_im_out(792)
        );

 
    UMUL_793 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(793),
            data_im_in => first_stage_im_out(793),
            re_multiplicator => "0010011011000001", --- 0.605529785156 + j-0.795837402344
            im_multiplicator => "1100110100010001",
            data_re_out => mul_re_out(793),
            data_im_out => mul_im_out(793)
        );

 
    UMUL_794 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(794),
            data_im_in => first_stage_im_out(794),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j-0.817565917969
            im_multiplicator => "1100101110101101",
            data_re_out => mul_re_out(794),
            data_im_out => mul_im_out(794)
        );

 
    UMUL_795 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(795),
            data_im_in => first_stage_im_out(795),
            re_multiplicator => "0010001011100111", --- 0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(795),
            data_im_out => mul_im_out(795)
        );

 
    UMUL_796 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(796),
            data_im_in => first_stage_im_out(796),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(796),
            data_im_out => mul_im_out(796)
        );

 
    UMUL_797 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(797),
            data_im_in => first_stage_im_out(797),
            re_multiplicator => "0001111011011100", --- 0.482177734375 + j-0.876098632812
            im_multiplicator => "1100011111101110",
            data_re_out => mul_re_out(797),
            data_im_out => mul_im_out(797)
        );

 
    UMUL_798 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(798),
            data_im_in => first_stage_im_out(798),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(798),
            data_im_out => mul_im_out(798)
        );

 
    UMUL_799 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(799),
            data_im_in => first_stage_im_out(799),
            re_multiplicator => "0001101010100111", --- 0.416442871094 + j-0.9091796875
            im_multiplicator => "1100010111010000",
            data_re_out => mul_re_out(799),
            data_im_out => mul_im_out(799)
        );

 
    UMUL_800 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(800),
            data_im_in => first_stage_im_out(800),
            re_multiplicator => "0001100001111110", --- 0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(800),
            data_im_out => mul_im_out(800)
        );

 
    UMUL_801 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(801),
            data_im_in => first_stage_im_out(801),
            re_multiplicator => "0001011001001100", --- 0.348388671875 + j-0.937316894531
            im_multiplicator => "1100010000000011",
            data_re_out => mul_re_out(801),
            data_im_out => mul_im_out(801)
        );

 
    UMUL_802 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(802),
            data_im_in => first_stage_im_out(802),
            re_multiplicator => "0001010000010011", --- 0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(802),
            data_im_out => mul_im_out(802)
        );

 
    UMUL_803 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(803),
            data_im_in => first_stage_im_out(803),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(803),
            data_im_out => mul_im_out(803)
        );

 
    UMUL_804 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(804),
            data_im_in => first_stage_im_out(804),
            re_multiplicator => "0000111110001101", --- 0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(804),
            data_im_out => mul_im_out(804)
        );

 
    UMUL_805 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(805),
            data_im_in => first_stage_im_out(805),
            re_multiplicator => "0000110101000001", --- 0.207092285156 + j-0.978332519531
            im_multiplicator => "1100000101100011",
            data_re_out => mul_re_out(805),
            data_im_out => mul_im_out(805)
        );

 
    UMUL_806 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(806),
            data_im_in => first_stage_im_out(806),
            re_multiplicator => "0000101011110001", --- 0.170959472656 + j-0.985290527344
            im_multiplicator => "1100000011110001",
            data_re_out => mul_re_out(806),
            data_im_out => mul_im_out(806)
        );

 
    UMUL_807 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(807),
            data_im_in => first_stage_im_out(807),
            re_multiplicator => "0000100010011101", --- 0.134582519531 + j-0.990905761719
            im_multiplicator => "1100000010010101",
            data_re_out => mul_re_out(807),
            data_im_out => mul_im_out(807)
        );

 
    UMUL_808 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(808),
            data_im_in => first_stage_im_out(808),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(808),
            data_im_out => mul_im_out(808)
        );

 
    UMUL_809 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(809),
            data_im_in => first_stage_im_out(809),
            re_multiplicator => "0000001111101101", --- 0.0613403320312 + j-0.998107910156
            im_multiplicator => "1100000000011111",
            data_re_out => mul_re_out(809),
            data_im_out => mul_im_out(809)
        );

 
    UMUL_810 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(810),
            data_im_in => first_stage_im_out(810),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(810),
            data_im_out => mul_im_out(810)
        );

 
    UMUL_811 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(811),
            data_im_in => first_stage_im_out(811),
            re_multiplicator => "1111111100110111", --- -0.0122680664062 + j-0.999938964844
            im_multiplicator => "1100000000000001",
            data_re_out => mul_re_out(811),
            data_im_out => mul_im_out(811)
        );

 
    UMUL_812 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(812),
            data_im_in => first_stage_im_out(812),
            re_multiplicator => "1111110011011100", --- -0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(812),
            data_im_out => mul_im_out(812)
        );

 
    UMUL_813 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(813),
            data_im_in => first_stage_im_out(813),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(813),
            data_im_out => mul_im_out(813)
        );

 
    UMUL_814 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(814),
            data_im_in => first_stage_im_out(814),
            re_multiplicator => "1111100000101010", --- -0.122436523438 + j-0.992492675781
            im_multiplicator => "1100000001111011",
            data_re_out => mul_re_out(814),
            data_im_out => mul_im_out(814)
        );

 
    UMUL_815 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(815),
            data_im_in => first_stage_im_out(815),
            re_multiplicator => "1111010111010101", --- -0.158874511719 + j-0.9873046875
            im_multiplicator => "1100000011010000",
            data_re_out => mul_re_out(815),
            data_im_out => mul_im_out(815)
        );

 
    UMUL_816 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(816),
            data_im_in => first_stage_im_out(816),
            re_multiplicator => "1111001110000100", --- -0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(816),
            data_im_out => mul_im_out(816)
        );

 
    UMUL_817 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(817),
            data_im_in => first_stage_im_out(817),
            re_multiplicator => "1111000100110110", --- -0.231079101562 + j-0.972961425781
            im_multiplicator => "1100000110111011",
            data_re_out => mul_re_out(817),
            data_im_out => mul_im_out(817)
        );

 
    UMUL_818 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(818),
            data_im_in => first_stage_im_out(818),
            re_multiplicator => "1110111011101110", --- -0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(818),
            data_im_out => mul_im_out(818)
        );

 
    UMUL_819 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(819),
            data_im_in => first_stage_im_out(819),
            re_multiplicator => "1110110010101100", --- -0.302001953125 + j-0.953308105469
            im_multiplicator => "1100001011111101",
            data_re_out => mul_re_out(819),
            data_im_out => mul_im_out(819)
        );

 
    UMUL_820 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(820),
            data_im_in => first_stage_im_out(820),
            re_multiplicator => "1110101001110000", --- -0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(820),
            data_im_out => mul_im_out(820)
        );

 
    UMUL_821 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(821),
            data_im_in => first_stage_im_out(821),
            re_multiplicator => "1110100000111100", --- -0.371337890625 + j-0.928527832031
            im_multiplicator => "1100010010010011",
            data_re_out => mul_re_out(821),
            data_im_out => mul_im_out(821)
        );

 
    UMUL_822 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(822),
            data_im_in => first_stage_im_out(822),
            re_multiplicator => "1110011000010001", --- -0.405212402344 + j-0.914184570312
            im_multiplicator => "1100010101111110",
            data_re_out => mul_re_out(822),
            data_im_out => mul_im_out(822)
        );

 
    UMUL_823 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(823),
            data_im_in => first_stage_im_out(823),
            re_multiplicator => "1110001111101110", --- -0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(823),
            data_im_out => mul_im_out(823)
        );

 
    UMUL_824 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(824),
            data_im_in => first_stage_im_out(824),
            re_multiplicator => "1110000111010101", --- -0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(824),
            data_im_out => mul_im_out(824)
        );

 
    UMUL_825 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(825),
            data_im_in => first_stage_im_out(825),
            re_multiplicator => "1101111111000110", --- -0.503540039062 + j-0.863952636719
            im_multiplicator => "1100100010110101",
            data_re_out => mul_re_out(825),
            data_im_out => mul_im_out(825)
        );

 
    UMUL_826 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(826),
            data_im_in => first_stage_im_out(826),
            re_multiplicator => "1101110111000011", --- -0.534973144531 + j-0.844848632812
            im_multiplicator => "1100100111101110",
            data_re_out => mul_re_out(826),
            data_im_out => mul_im_out(826)
        );

 
    UMUL_827 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(827),
            data_im_in => first_stage_im_out(827),
            re_multiplicator => "1101101111001011", --- -0.565734863281 + j-0.824584960938
            im_multiplicator => "1100101100111010",
            data_re_out => mul_re_out(827),
            data_im_out => mul_im_out(827)
        );

 
    UMUL_828 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(828),
            data_im_in => first_stage_im_out(828),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(828),
            data_im_out => mul_im_out(828)
        );

 
    UMUL_829 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(829),
            data_im_in => first_stage_im_out(829),
            re_multiplicator => "1101100000000010", --- -0.624877929688 + j-0.78076171875
            im_multiplicator => "1100111000001000",
            data_re_out => mul_re_out(829),
            data_im_out => mul_im_out(829)
        );

 
    UMUL_830 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(830),
            data_im_in => first_stage_im_out(830),
            re_multiplicator => "1101011000110010", --- -0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(830),
            data_im_out => mul_im_out(830)
        );

 
    UMUL_831 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(831),
            data_im_in => first_stage_im_out(831),
            re_multiplicator => "1101010001110001", --- -0.680603027344 + j-0.732666015625
            im_multiplicator => "1101000100011100",
            data_re_out => mul_re_out(831),
            data_im_out => mul_im_out(831)
        );

 
    UMUL_832 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(832),
            data_im_in => first_stage_im_out(832),
            data_re_out => mul_re_out(832),
            data_im_out => mul_im_out(832)
        );

 
    UMUL_833 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(833),
            data_im_in => first_stage_im_out(833),
            re_multiplicator => "0011111111110011", --- 0.999206542969 + j-0.0398559570312
            im_multiplicator => "1111110101110011",
            data_re_out => mul_re_out(833),
            data_im_out => mul_im_out(833)
        );

 
    UMUL_834 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(834),
            data_im_in => first_stage_im_out(834),
            re_multiplicator => "0011111111001100", --- 0.996826171875 + j-0.0797119140625
            im_multiplicator => "1111101011100110",
            data_re_out => mul_re_out(834),
            data_im_out => mul_im_out(834)
        );

 
    UMUL_835 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(835),
            data_im_in => first_stage_im_out(835),
            re_multiplicator => "0011111110001011", --- 0.992858886719 + j-0.119384765625
            im_multiplicator => "1111100001011100",
            data_re_out => mul_re_out(835),
            data_im_out => mul_im_out(835)
        );

 
    UMUL_836 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(836),
            data_im_in => first_stage_im_out(836),
            re_multiplicator => "0011111100110000", --- 0.9873046875 + j-0.158874511719
            im_multiplicator => "1111010111010101",
            data_re_out => mul_re_out(836),
            data_im_out => mul_im_out(836)
        );

 
    UMUL_837 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(837),
            data_im_in => first_stage_im_out(837),
            re_multiplicator => "0011111010111011", --- 0.980163574219 + j-0.198120117188
            im_multiplicator => "1111001101010010",
            data_re_out => mul_re_out(837),
            data_im_out => mul_im_out(837)
        );

 
    UMUL_838 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(838),
            data_im_in => first_stage_im_out(838),
            re_multiplicator => "0011111000101101", --- 0.971496582031 + j-0.236999511719
            im_multiplicator => "1111000011010101",
            data_re_out => mul_re_out(838),
            data_im_out => mul_im_out(838)
        );

 
    UMUL_839 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(839),
            data_im_in => first_stage_im_out(839),
            re_multiplicator => "0011110110000110", --- 0.961303710938 + j-0.275573730469
            im_multiplicator => "1110111001011101",
            data_re_out => mul_re_out(839),
            data_im_out => mul_im_out(839)
        );

 
    UMUL_840 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(840),
            data_im_in => first_stage_im_out(840),
            re_multiplicator => "0011110011000101", --- 0.949523925781 + j-0.313659667969
            im_multiplicator => "1110101111101101",
            data_re_out => mul_re_out(840),
            data_im_out => mul_im_out(840)
        );

 
    UMUL_841 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(841),
            data_im_in => first_stage_im_out(841),
            re_multiplicator => "0011101111101100", --- 0.936279296875 + j-0.351318359375
            im_multiplicator => "1110100110000100",
            data_re_out => mul_re_out(841),
            data_im_out => mul_im_out(841)
        );

 
    UMUL_842 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(842),
            data_im_in => first_stage_im_out(842),
            re_multiplicator => "0011101011111010", --- 0.921508789062 + j-0.388366699219
            im_multiplicator => "1110011100100101",
            data_re_out => mul_re_out(842),
            data_im_out => mul_im_out(842)
        );

 
    UMUL_843 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(843),
            data_im_in => first_stage_im_out(843),
            re_multiplicator => "0011100111110000", --- 0.9052734375 + j-0.4248046875
            im_multiplicator => "1110010011010000",
            data_re_out => mul_re_out(843),
            data_im_out => mul_im_out(843)
        );

 
    UMUL_844 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(844),
            data_im_in => first_stage_im_out(844),
            re_multiplicator => "0011100011001111", --- 0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(844),
            data_im_out => mul_im_out(844)
        );

 
    UMUL_845 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(845),
            data_im_in => first_stage_im_out(845),
            re_multiplicator => "0011011110010111", --- 0.868591308594 + j-0.495544433594
            im_multiplicator => "1110000001001001",
            data_re_out => mul_re_out(845),
            data_im_out => mul_im_out(845)
        );

 
    UMUL_846 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(846),
            data_im_in => first_stage_im_out(846),
            re_multiplicator => "0011011001001000", --- 0.84814453125 + j-0.52978515625
            im_multiplicator => "1101111000011000",
            data_re_out => mul_re_out(846),
            data_im_out => mul_im_out(846)
        );

 
    UMUL_847 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(847),
            data_im_in => first_stage_im_out(847),
            re_multiplicator => "0011010011100010", --- 0.826293945312 + j-0.563171386719
            im_multiplicator => "1101101111110101",
            data_re_out => mul_re_out(847),
            data_im_out => mul_im_out(847)
        );

 
    UMUL_848 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(848),
            data_im_in => first_stage_im_out(848),
            re_multiplicator => "0011001101101000", --- 0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(848),
            data_im_out => mul_im_out(848)
        );

 
    UMUL_849 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(849),
            data_im_in => first_stage_im_out(849),
            re_multiplicator => "0011000111011000", --- 0.77880859375 + j-0.627258300781
            im_multiplicator => "1101011111011011",
            data_re_out => mul_re_out(849),
            data_im_out => mul_im_out(849)
        );

 
    UMUL_850 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(850),
            data_im_in => first_stage_im_out(850),
            re_multiplicator => "0011000000110100", --- 0.753173828125 + j-0.657836914062
            im_multiplicator => "1101010111100110",
            data_re_out => mul_re_out(850),
            data_im_out => mul_im_out(850)
        );

 
    UMUL_851 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(851),
            data_im_in => first_stage_im_out(851),
            re_multiplicator => "0010111001111101", --- 0.726379394531 + j-0.687316894531
            im_multiplicator => "1101010000000011",
            data_re_out => mul_re_out(851),
            data_im_out => mul_im_out(851)
        );

 
    UMUL_852 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(852),
            data_im_in => first_stage_im_out(852),
            re_multiplicator => "0010110010110010", --- 0.698364257812 + j-0.715759277344
            im_multiplicator => "1101001000110001",
            data_re_out => mul_re_out(852),
            data_im_out => mul_im_out(852)
        );

 
    UMUL_853 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(853),
            data_im_in => first_stage_im_out(853),
            re_multiplicator => "0010101011010110", --- 0.669311523438 + j-0.742980957031
            im_multiplicator => "1101000001110011",
            data_re_out => mul_re_out(853),
            data_im_out => mul_im_out(853)
        );

 
    UMUL_854 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(854),
            data_im_in => first_stage_im_out(854),
            re_multiplicator => "0010100011100111", --- 0.639099121094 + j-0.769104003906
            im_multiplicator => "1100111011000111",
            data_re_out => mul_re_out(854),
            data_im_out => mul_im_out(854)
        );

 
    UMUL_855 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(855),
            data_im_in => first_stage_im_out(855),
            re_multiplicator => "0010011011101001", --- 0.607971191406 + j-0.7939453125
            im_multiplicator => "1100110100110000",
            data_re_out => mul_re_out(855),
            data_im_out => mul_im_out(855)
        );

 
    UMUL_856 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(856),
            data_im_in => first_stage_im_out(856),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j-0.817565917969
            im_multiplicator => "1100101110101101",
            data_re_out => mul_re_out(856),
            data_im_out => mul_im_out(856)
        );

 
    UMUL_857 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(857),
            data_im_in => first_stage_im_out(857),
            re_multiplicator => "0010001010111100", --- 0.542724609375 + j-0.839904785156
            im_multiplicator => "1100101000111111",
            data_re_out => mul_re_out(857),
            data_im_out => mul_im_out(857)
        );

 
    UMUL_858 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(858),
            data_im_in => first_stage_im_out(858),
            re_multiplicator => "0010000010010001", --- 0.508850097656 + j-0.86083984375
            im_multiplicator => "1100100011101000",
            data_re_out => mul_re_out(858),
            data_im_out => mul_im_out(858)
        );

 
    UMUL_859 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(859),
            data_im_in => first_stage_im_out(859),
            re_multiplicator => "0001111001011000", --- 0.47412109375 + j-0.880493164062
            im_multiplicator => "1100011110100110",
            data_re_out => mul_re_out(859),
            data_im_out => mul_im_out(859)
        );

 
    UMUL_860 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(860),
            data_im_in => first_stage_im_out(860),
            re_multiplicator => "0001110000010010", --- 0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(860),
            data_im_out => mul_im_out(860)
        );

 
    UMUL_861 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(861),
            data_im_in => first_stage_im_out(861),
            re_multiplicator => "0001100111000001", --- 0.402404785156 + j-0.915466308594
            im_multiplicator => "1100010101101001",
            data_re_out => mul_re_out(861),
            data_im_out => mul_im_out(861)
        );

 
    UMUL_862 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(862),
            data_im_in => first_stage_im_out(862),
            re_multiplicator => "0001011101100110", --- 0.365600585938 + j-0.930786132812
            im_multiplicator => "1100010001101110",
            data_re_out => mul_re_out(862),
            data_im_out => mul_im_out(862)
        );

 
    UMUL_863 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(863),
            data_im_in => first_stage_im_out(863),
            re_multiplicator => "0001010100000001", --- 0.328186035156 + j-0.944580078125
            im_multiplicator => "1100001110001100",
            data_re_out => mul_re_out(863),
            data_im_out => mul_im_out(863)
        );

 
    UMUL_864 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(864),
            data_im_in => first_stage_im_out(864),
            re_multiplicator => "0001001010010100", --- 0.290283203125 + j-0.956970214844
            im_multiplicator => "1100001011000001",
            data_re_out => mul_re_out(864),
            data_im_out => mul_im_out(864)
        );

 
    UMUL_865 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(865),
            data_im_in => first_stage_im_out(865),
            re_multiplicator => "0001000000011111", --- 0.251892089844 + j-0.9677734375
            im_multiplicator => "1100001000010000",
            data_re_out => mul_re_out(865),
            data_im_out => mul_im_out(865)
        );

 
    UMUL_866 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(866),
            data_im_in => first_stage_im_out(866),
            re_multiplicator => "0000110110100100", --- 0.213134765625 + j-0.97705078125
            im_multiplicator => "1100000101111000",
            data_re_out => mul_re_out(866),
            data_im_out => mul_im_out(866)
        );

 
    UMUL_867 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(867),
            data_im_in => first_stage_im_out(867),
            re_multiplicator => "0000101100100011", --- 0.174011230469 + j-0.984741210938
            im_multiplicator => "1100000011111010",
            data_re_out => mul_re_out(867),
            data_im_out => mul_im_out(867)
        );

 
    UMUL_868 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(868),
            data_im_in => first_stage_im_out(868),
            re_multiplicator => "0000100010011101", --- 0.134582519531 + j-0.990905761719
            im_multiplicator => "1100000010010101",
            data_re_out => mul_re_out(868),
            data_im_out => mul_im_out(868)
        );

 
    UMUL_869 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(869),
            data_im_in => first_stage_im_out(869),
            re_multiplicator => "0000011000010100", --- 0.094970703125 + j-0.995483398438
            im_multiplicator => "1100000001001010",
            data_re_out => mul_re_out(869),
            data_im_out => mul_im_out(869)
        );

 
    UMUL_870 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(870),
            data_im_in => first_stage_im_out(870),
            re_multiplicator => "0000001110001000", --- 0.05517578125 + j-0.998474121094
            im_multiplicator => "1100000000011001",
            data_re_out => mul_re_out(870),
            data_im_out => mul_im_out(870)
        );

 
    UMUL_871 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(871),
            data_im_in => first_stage_im_out(871),
            re_multiplicator => "0000000011111011", --- 0.0153198242188 + j-0.999877929688
            im_multiplicator => "1100000000000010",
            data_re_out => mul_re_out(871),
            data_im_out => mul_im_out(871)
        );

 
    UMUL_872 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(872),
            data_im_in => first_stage_im_out(872),
            re_multiplicator => "1111111001101110", --- -0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(872),
            data_im_out => mul_im_out(872)
        );

 
    UMUL_873 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(873),
            data_im_in => first_stage_im_out(873),
            re_multiplicator => "1111101111100001", --- -0.0643920898438 + j-0.997924804688
            im_multiplicator => "1100000000100010",
            data_re_out => mul_re_out(873),
            data_im_out => mul_im_out(873)
        );

 
    UMUL_874 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(874),
            data_im_in => first_stage_im_out(874),
            re_multiplicator => "1111100101010110", --- -0.104125976562 + j-0.994567871094
            im_multiplicator => "1100000001011001",
            data_re_out => mul_re_out(874),
            data_im_out => mul_im_out(874)
        );

 
    UMUL_875 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(875),
            data_im_in => first_stage_im_out(875),
            re_multiplicator => "1111011011001110", --- -0.143676757812 + j-0.989624023438
            im_multiplicator => "1100000010101010",
            data_re_out => mul_re_out(875),
            data_im_out => mul_im_out(875)
        );

 
    UMUL_876 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(876),
            data_im_in => first_stage_im_out(876),
            re_multiplicator => "1111010001001001", --- -0.183044433594 + j-0.983093261719
            im_multiplicator => "1100000100010101",
            data_re_out => mul_re_out(876),
            data_im_out => mul_im_out(876)
        );

 
    UMUL_877 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(877),
            data_im_in => first_stage_im_out(877),
            re_multiplicator => "1111000111001001", --- -0.222106933594 + j-0.975036621094
            im_multiplicator => "1100000110011001",
            data_re_out => mul_re_out(877),
            data_im_out => mul_im_out(877)
        );

 
    UMUL_878 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(878),
            data_im_in => first_stage_im_out(878),
            re_multiplicator => "1110111101001111", --- -0.260803222656 + j-0.965393066406
            im_multiplicator => "1100001000110111",
            data_re_out => mul_re_out(878),
            data_im_out => mul_im_out(878)
        );

 
    UMUL_879 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(879),
            data_im_in => first_stage_im_out(879),
            re_multiplicator => "1110110011011100", --- -0.299072265625 + j-0.954223632812
            im_multiplicator => "1100001011101110",
            data_re_out => mul_re_out(879),
            data_im_out => mul_im_out(879)
        );

 
    UMUL_880 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(880),
            data_im_in => first_stage_im_out(880),
            re_multiplicator => "1110101001110000", --- -0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(880),
            data_im_out => mul_im_out(880)
        );

 
    UMUL_881 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(881),
            data_im_in => first_stage_im_out(881),
            re_multiplicator => "1110100000001110", --- -0.374145507812 + j-0.927368164062
            im_multiplicator => "1100010010100110",
            data_re_out => mul_re_out(881),
            data_im_out => mul_im_out(881)
        );

 
    UMUL_882 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(882),
            data_im_in => first_stage_im_out(882),
            re_multiplicator => "1110010110110101", --- -0.410827636719 + j-0.911682128906
            im_multiplicator => "1100010110100111",
            data_re_out => mul_re_out(882),
            data_im_out => mul_im_out(882)
        );

 
    UMUL_883 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(883),
            data_im_in => first_stage_im_out(883),
            re_multiplicator => "1110001101100111", --- -0.446838378906 + j-0.894592285156
            im_multiplicator => "1100011010111111",
            data_re_out => mul_re_out(883),
            data_im_out => mul_im_out(883)
        );

 
    UMUL_884 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(884),
            data_im_in => first_stage_im_out(884),
            re_multiplicator => "1110000100100100", --- -0.482177734375 + j-0.876098632812
            im_multiplicator => "1100011111101110",
            data_re_out => mul_re_out(884),
            data_im_out => mul_im_out(884)
        );

 
    UMUL_885 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(885),
            data_im_in => first_stage_im_out(885),
            re_multiplicator => "1101111011101110", --- -0.516723632812 + j-0.856140136719
            im_multiplicator => "1100100100110101",
            data_re_out => mul_re_out(885),
            data_im_out => mul_im_out(885)
        );

 
    UMUL_886 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(886),
            data_im_in => first_stage_im_out(886),
            re_multiplicator => "1101110011000101", --- -0.550476074219 + j-0.834838867188
            im_multiplicator => "1100101010010010",
            data_re_out => mul_re_out(886),
            data_im_out => mul_im_out(886)
        );

 
    UMUL_887 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(887),
            data_im_in => first_stage_im_out(887),
            re_multiplicator => "1101101010101011", --- -0.583312988281 + j-0.812255859375
            im_multiplicator => "1100110000000100",
            data_re_out => mul_re_out(887),
            data_im_out => mul_im_out(887)
        );

 
    UMUL_888 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(888),
            data_im_in => first_stage_im_out(888),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j-0.788330078125
            im_multiplicator => "1100110110001100",
            data_re_out => mul_re_out(888),
            data_im_out => mul_im_out(888)
        );

 
    UMUL_889 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(889),
            data_im_in => first_stage_im_out(889),
            re_multiplicator => "1101011010100101", --- -0.646179199219 + j-0.76318359375
            im_multiplicator => "1100111100101000",
            data_re_out => mul_re_out(889),
            data_im_out => mul_im_out(889)
        );

 
    UMUL_890 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(890),
            data_im_in => first_stage_im_out(890),
            re_multiplicator => "1101010010111011", --- -0.676086425781 + j-0.73681640625
            im_multiplicator => "1101000011011000",
            data_re_out => mul_re_out(890),
            data_im_out => mul_im_out(890)
        );

 
    UMUL_891 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(891),
            data_im_in => first_stage_im_out(891),
            re_multiplicator => "1101001011100010", --- -0.704956054688 + j-0.709289550781
            im_multiplicator => "1101001010011011",
            data_re_out => mul_re_out(891),
            data_im_out => mul_im_out(891)
        );

 
    UMUL_892 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(892),
            data_im_in => first_stage_im_out(892),
            re_multiplicator => "1101000100011100", --- -0.732666015625 + j-0.680603027344
            im_multiplicator => "1101010001110001",
            data_re_out => mul_re_out(892),
            data_im_out => mul_im_out(892)
        );

 
    UMUL_893 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(893),
            data_im_in => first_stage_im_out(893),
            re_multiplicator => "1100111101101001", --- -0.759216308594 + j-0.650817871094
            im_multiplicator => "1101011001011001",
            data_re_out => mul_re_out(893),
            data_im_out => mul_im_out(893)
        );

 
    UMUL_894 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(894),
            data_im_in => first_stage_im_out(894),
            re_multiplicator => "1100110111001010", --- -0.784545898438 + j-0.620056152344
            im_multiplicator => "1101100001010001",
            data_re_out => mul_re_out(894),
            data_im_out => mul_im_out(894)
        );

 
    UMUL_895 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(895),
            data_im_in => first_stage_im_out(895),
            re_multiplicator => "1100110000111111", --- -0.808654785156 + j-0.588256835938
            im_multiplicator => "1101101001011010",
            data_re_out => mul_re_out(895),
            data_im_out => mul_im_out(895)
        );

 
    UMUL_896 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(896),
            data_im_in => first_stage_im_out(896),
            data_re_out => mul_re_out(896),
            data_im_out => mul_im_out(896)
        );

 
    UMUL_897 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(897),
            data_im_in => first_stage_im_out(897),
            re_multiplicator => "0011111111110001", --- 0.999084472656 + j-0.04296875
            im_multiplicator => "1111110101000000",
            data_re_out => mul_re_out(897),
            data_im_out => mul_im_out(897)
        );

 
    UMUL_898 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(898),
            data_im_in => first_stage_im_out(898),
            re_multiplicator => "0011111111000100", --- 0.996337890625 + j-0.0858154296875
            im_multiplicator => "1111101010000010",
            data_re_out => mul_re_out(898),
            data_im_out => mul_im_out(898)
        );

 
    UMUL_899 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(899),
            data_im_in => first_stage_im_out(899),
            re_multiplicator => "0011111101111000", --- 0.99169921875 + j-0.128479003906
            im_multiplicator => "1111011111000111",
            data_re_out => mul_re_out(899),
            data_im_out => mul_im_out(899)
        );

 
    UMUL_900 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(900),
            data_im_in => first_stage_im_out(900),
            re_multiplicator => "0011111100001111", --- 0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(900),
            data_im_out => mul_im_out(900)
        );

 
    UMUL_901 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(901),
            data_im_in => first_stage_im_out(901),
            re_multiplicator => "0011111010001000", --- 0.97705078125 + j-0.213134765625
            im_multiplicator => "1111001001011100",
            data_re_out => mul_re_out(901),
            data_im_out => mul_im_out(901)
        );

 
    UMUL_902 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(902),
            data_im_in => first_stage_im_out(902),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(902),
            data_im_out => mul_im_out(902)
        );

 
    UMUL_903 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(903),
            data_im_in => first_stage_im_out(903),
            re_multiplicator => "0011110100100001", --- 0.955139160156 + j-0.296142578125
            im_multiplicator => "1110110100001100",
            data_re_out => mul_re_out(903),
            data_im_out => mul_im_out(903)
        );

 
    UMUL_904 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(904),
            data_im_in => first_stage_im_out(904),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(904),
            data_im_out => mul_im_out(904)
        );

 
    UMUL_905 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(905),
            data_im_in => first_stage_im_out(905),
            re_multiplicator => "0011101101000111", --- 0.926208496094 + j-0.377014160156
            im_multiplicator => "1110011111011111",
            data_re_out => mul_re_out(905),
            data_im_out => mul_im_out(905)
        );

 
    UMUL_906 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(906),
            data_im_in => first_stage_im_out(906),
            re_multiplicator => "0011101000110000", --- 0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(906),
            data_im_out => mul_im_out(906)
        );

 
    UMUL_907 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(907),
            data_im_in => first_stage_im_out(907),
            re_multiplicator => "0011100011111101", --- 0.890441894531 + j-0.455078125
            im_multiplicator => "1110001011100000",
            data_re_out => mul_re_out(907),
            data_im_out => mul_im_out(907)
        );

 
    UMUL_908 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(908),
            data_im_in => first_stage_im_out(908),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(908),
            data_im_out => mul_im_out(908)
        );

 
    UMUL_909 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(909),
            data_im_in => first_stage_im_out(909),
            re_multiplicator => "0011011001001000", --- 0.84814453125 + j-0.52978515625
            im_multiplicator => "1101111000011000",
            data_re_out => mul_re_out(909),
            data_im_out => mul_im_out(909)
        );

 
    UMUL_910 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(910),
            data_im_in => first_stage_im_out(910),
            re_multiplicator => "0011010011000110", --- 0.824584960938 + j-0.565734863281
            im_multiplicator => "1101101111001011",
            data_re_out => mul_re_out(910),
            data_im_out => mul_im_out(910)
        );

 
    UMUL_911 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(911),
            data_im_in => first_stage_im_out(911),
            re_multiplicator => "0011001100101100", --- 0.799560546875 + j-0.600646972656
            im_multiplicator => "1101100110001111",
            data_re_out => mul_re_out(911),
            data_im_out => mul_im_out(911)
        );

 
    UMUL_912 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(912),
            data_im_in => first_stage_im_out(912),
            re_multiplicator => "0011000101111001", --- 0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(912),
            data_im_out => mul_im_out(912)
        );

 
    UMUL_913 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(913),
            data_im_in => first_stage_im_out(913),
            re_multiplicator => "0010111110101111", --- 0.745056152344 + j-0.6669921875
            im_multiplicator => "1101010101010000",
            data_re_out => mul_re_out(913),
            data_im_out => mul_im_out(913)
        );

 
    UMUL_914 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(914),
            data_im_in => first_stage_im_out(914),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(914),
            data_im_out => mul_im_out(914)
        );

 
    UMUL_915 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(915),
            data_im_in => first_stage_im_out(915),
            re_multiplicator => "0010101111011000", --- 0.68505859375 + j-0.728454589844
            im_multiplicator => "1101000101100001",
            data_re_out => mul_re_out(915),
            data_im_out => mul_im_out(915)
        );

 
    UMUL_916 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(916),
            data_im_in => first_stage_im_out(916),
            re_multiplicator => "0010100111001110", --- 0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(916),
            data_im_out => mul_im_out(916)
        );

 
    UMUL_917 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(917),
            data_im_in => first_stage_im_out(917),
            re_multiplicator => "0010011110101111", --- 0.620056152344 + j-0.784545898438
            im_multiplicator => "1100110111001010",
            data_re_out => mul_re_out(917),
            data_im_out => mul_im_out(917)
        );

 
    UMUL_918 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(918),
            data_im_in => first_stage_im_out(918),
            re_multiplicator => "0010010101111110", --- 0.585815429688 + j-0.810485839844
            im_multiplicator => "1100110000100001",
            data_re_out => mul_re_out(918),
            data_im_out => mul_im_out(918)
        );

 
    UMUL_919 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(919),
            data_im_in => first_stage_im_out(919),
            re_multiplicator => "0010001100111011", --- 0.550476074219 + j-0.834838867188
            im_multiplicator => "1100101010010010",
            data_re_out => mul_re_out(919),
            data_im_out => mul_im_out(919)
        );

 
    UMUL_920 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(920),
            data_im_in => first_stage_im_out(920),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(920),
            data_im_out => mul_im_out(920)
        );

 
    UMUL_921 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(921),
            data_im_in => first_stage_im_out(921),
            re_multiplicator => "0001111010000100", --- 0.476806640625 + j-0.879028320312
            im_multiplicator => "1100011110111110",
            data_re_out => mul_re_out(921),
            data_im_out => mul_im_out(921)
        );

 
    UMUL_922 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(922),
            data_im_in => first_stage_im_out(922),
            re_multiplicator => "0001110000010010", --- 0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(922),
            data_im_out => mul_im_out(922)
        );

 
    UMUL_923 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(923),
            data_im_in => first_stage_im_out(923),
            re_multiplicator => "0001100110010011", --- 0.399597167969 + j-0.916687011719
            im_multiplicator => "1100010101010101",
            data_re_out => mul_re_out(923),
            data_im_out => mul_im_out(923)
        );

 
    UMUL_924 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(924),
            data_im_in => first_stage_im_out(924),
            re_multiplicator => "0001011100001001", --- 0.359924316406 + j-0.932983398438
            im_multiplicator => "1100010001001010",
            data_re_out => mul_re_out(924),
            data_im_out => mul_im_out(924)
        );

 
    UMUL_925 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(925),
            data_im_in => first_stage_im_out(925),
            re_multiplicator => "0001010001110011", --- 0.319519042969 + j-0.947570800781
            im_multiplicator => "1100001101011011",
            data_re_out => mul_re_out(925),
            data_im_out => mul_im_out(925)
        );

 
    UMUL_926 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(926),
            data_im_in => first_stage_im_out(926),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(926),
            data_im_out => mul_im_out(926)
        );

 
    UMUL_927 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(927),
            data_im_in => first_stage_im_out(927),
            re_multiplicator => "0000111100101011", --- 0.236999511719 + j-0.971496582031
            im_multiplicator => "1100000111010011",
            data_re_out => mul_re_out(927),
            data_im_out => mul_im_out(927)
        );

 
    UMUL_928 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(928),
            data_im_in => first_stage_im_out(928),
            re_multiplicator => "0000110001111100", --- 0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(928),
            data_im_out => mul_im_out(928)
        );

 
    UMUL_929 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(929),
            data_im_in => first_stage_im_out(929),
            re_multiplicator => "0000100111000111", --- 0.152770996094 + j-0.98828125
            im_multiplicator => "1100000011000000",
            data_re_out => mul_re_out(929),
            data_im_out => mul_im_out(929)
        );

 
    UMUL_930 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(930),
            data_im_in => first_stage_im_out(930),
            re_multiplicator => "0000011100001110", --- 0.110229492188 + j-0.993896484375
            im_multiplicator => "1100000001100100",
            data_re_out => mul_re_out(930),
            data_im_out => mul_im_out(930)
        );

 
    UMUL_931 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(931),
            data_im_in => first_stage_im_out(931),
            re_multiplicator => "0000010001010001", --- 0.0674438476562 + j-0.997741699219
            im_multiplicator => "1100000000100101",
            data_re_out => mul_re_out(931),
            data_im_out => mul_im_out(931)
        );

 
    UMUL_932 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(932),
            data_im_in => first_stage_im_out(932),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(932),
            data_im_out => mul_im_out(932)
        );

 
    UMUL_933 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(933),
            data_im_in => first_stage_im_out(933),
            re_multiplicator => "1111111011010010", --- -0.0184326171875 + j-0.999816894531
            im_multiplicator => "1100000000000011",
            data_re_out => mul_re_out(933),
            data_im_out => mul_im_out(933)
        );

 
    UMUL_934 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(934),
            data_im_in => first_stage_im_out(934),
            re_multiplicator => "1111110000010011", --- -0.0613403320312 + j-0.998107910156
            im_multiplicator => "1100000000011111",
            data_re_out => mul_re_out(934),
            data_im_out => mul_im_out(934)
        );

 
    UMUL_935 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(935),
            data_im_in => first_stage_im_out(935),
            re_multiplicator => "1111100101010110", --- -0.104125976562 + j-0.994567871094
            im_multiplicator => "1100000001011001",
            data_re_out => mul_re_out(935),
            data_im_out => mul_im_out(935)
        );

 
    UMUL_936 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(936),
            data_im_in => first_stage_im_out(936),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(936),
            data_im_out => mul_im_out(936)
        );

 
    UMUL_937 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(937),
            data_im_in => first_stage_im_out(937),
            re_multiplicator => "1111001111100110", --- -0.189086914062 + j-0.98193359375
            im_multiplicator => "1100000100101000",
            data_re_out => mul_re_out(937),
            data_im_out => mul_im_out(937)
        );

 
    UMUL_938 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(938),
            data_im_in => first_stage_im_out(938),
            re_multiplicator => "1111000100110110", --- -0.231079101562 + j-0.972961425781
            im_multiplicator => "1100000110111011",
            data_re_out => mul_re_out(938),
            data_im_out => mul_im_out(938)
        );

 
    UMUL_939 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(939),
            data_im_in => first_stage_im_out(939),
            re_multiplicator => "1110111010001101", --- -0.272644042969 + j-0.962097167969
            im_multiplicator => "1100001001101101",
            data_re_out => mul_re_out(939),
            data_im_out => mul_im_out(939)
        );

 
    UMUL_940 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(940),
            data_im_in => first_stage_im_out(940),
            re_multiplicator => "1110101111101101", --- -0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(940),
            data_im_out => mul_im_out(940)
        );

 
    UMUL_941 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(941),
            data_im_in => first_stage_im_out(941),
            re_multiplicator => "1110100101010101", --- -0.354187011719 + j-0.935180664062
            im_multiplicator => "1100010000100110",
            data_re_out => mul_re_out(941),
            data_im_out => mul_im_out(941)
        );

 
    UMUL_942 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(942),
            data_im_in => first_stage_im_out(942),
            re_multiplicator => "1110011011001001", --- -0.393981933594 + j-0.919128417969
            im_multiplicator => "1100010100101101",
            data_re_out => mul_re_out(942),
            data_im_out => mul_im_out(942)
        );

 
    UMUL_943 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(943),
            data_im_in => first_stage_im_out(943),
            re_multiplicator => "1110010001001000", --- -0.43310546875 + j-0.9013671875
            im_multiplicator => "1100011001010000",
            data_re_out => mul_re_out(943),
            data_im_out => mul_im_out(943)
        );

 
    UMUL_944 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(944),
            data_im_in => first_stage_im_out(944),
            re_multiplicator => "1110000111010101", --- -0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(944),
            data_im_out => mul_im_out(944)
        );

 
    UMUL_945 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(945),
            data_im_in => first_stage_im_out(945),
            re_multiplicator => "1101111101101111", --- -0.508850097656 + j-0.86083984375
            im_multiplicator => "1100100011101000",
            data_re_out => mul_re_out(945),
            data_im_out => mul_im_out(945)
        );

 
    UMUL_946 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(946),
            data_im_in => first_stage_im_out(946),
            re_multiplicator => "1101110100011001", --- -0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(946),
            data_im_out => mul_im_out(946)
        );

 
    UMUL_947 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(947),
            data_im_in => first_stage_im_out(947),
            re_multiplicator => "1101101011010100", --- -0.580810546875 + j-0.814025878906
            im_multiplicator => "1100101111100111",
            data_re_out => mul_re_out(947),
            data_im_out => mul_im_out(947)
        );

 
    UMUL_948 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(948),
            data_im_in => first_stage_im_out(948),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j-0.788330078125
            im_multiplicator => "1100110110001100",
            data_re_out => mul_re_out(948),
            data_im_out => mul_im_out(948)
        );

 
    UMUL_949 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(949),
            data_im_in => first_stage_im_out(949),
            re_multiplicator => "1101011001111111", --- -0.648498535156 + j-0.76123046875
            im_multiplicator => "1100111101001000",
            data_re_out => mul_re_out(949),
            data_im_out => mul_im_out(949)
        );

 
    UMUL_950 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(950),
            data_im_in => first_stage_im_out(950),
            re_multiplicator => "1101010001110001", --- -0.680603027344 + j-0.732666015625
            im_multiplicator => "1101000100011100",
            data_re_out => mul_re_out(950),
            data_im_out => mul_im_out(950)
        );

 
    UMUL_951 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(951),
            data_im_in => first_stage_im_out(951),
            re_multiplicator => "1101001001111000", --- -0.71142578125 + j-0.702758789062
            im_multiplicator => "1101001100000110",
            data_re_out => mul_re_out(951),
            data_im_out => mul_im_out(951)
        );

 
    UMUL_952 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(952),
            data_im_in => first_stage_im_out(952),
            re_multiplicator => "1101000010010100", --- -0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(952),
            data_im_out => mul_im_out(952)
        );

 
    UMUL_953 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(953),
            data_im_in => first_stage_im_out(953),
            re_multiplicator => "1100111011000111", --- -0.769104003906 + j-0.639099121094
            im_multiplicator => "1101011100011001",
            data_re_out => mul_re_out(953),
            data_im_out => mul_im_out(953)
        );

 
    UMUL_954 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(954),
            data_im_in => first_stage_im_out(954),
            re_multiplicator => "1100110100010001", --- -0.795837402344 + j-0.605529785156
            im_multiplicator => "1101100100111111",
            data_re_out => mul_re_out(954),
            data_im_out => mul_im_out(954)
        );

 
    UMUL_955 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(955),
            data_im_in => first_stage_im_out(955),
            re_multiplicator => "1100101101110011", --- -0.821105957031 + j-0.57080078125
            im_multiplicator => "1101101101111000",
            data_re_out => mul_re_out(955),
            data_im_out => mul_im_out(955)
        );

 
    UMUL_956 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(956),
            data_im_in => first_stage_im_out(956),
            re_multiplicator => "1100100111101110", --- -0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(956),
            data_im_out => mul_im_out(956)
        );

 
    UMUL_957 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(957),
            data_im_in => first_stage_im_out(957),
            re_multiplicator => "1100100010000010", --- -0.867065429688 + j-0.498229980469
            im_multiplicator => "1110000000011101",
            data_re_out => mul_re_out(957),
            data_im_out => mul_im_out(957)
        );

 
    UMUL_958 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(958),
            data_im_in => first_stage_im_out(958),
            re_multiplicator => "1100011100110001", --- -0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(958),
            data_im_out => mul_im_out(958)
        );

 
    UMUL_959 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(959),
            data_im_in => first_stage_im_out(959),
            re_multiplicator => "1100010111111010", --- -0.906616210938 + j-0.421997070312
            im_multiplicator => "1110010011111110",
            data_re_out => mul_re_out(959),
            data_im_out => mul_im_out(959)
        );

 
    UMUL_960 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(960),
            data_im_in => first_stage_im_out(960),
            data_re_out => mul_re_out(960),
            data_im_out => mul_im_out(960)
        );

 
    UMUL_961 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(961),
            data_im_in => first_stage_im_out(961),
            re_multiplicator => "0011111111101111", --- 0.998962402344 + j-0.0460205078125
            im_multiplicator => "1111110100001110",
            data_re_out => mul_re_out(961),
            data_im_out => mul_im_out(961)
        );

 
    UMUL_962 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(962),
            data_im_in => first_stage_im_out(962),
            re_multiplicator => "0011111110111011", --- 0.995788574219 + j-0.0919189453125
            im_multiplicator => "1111101000011110",
            data_re_out => mul_re_out(962),
            data_im_out => mul_im_out(962)
        );

 
    UMUL_963 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(963),
            data_im_in => first_stage_im_out(963),
            re_multiplicator => "0011111101100100", --- 0.990478515625 + j-0.137634277344
            im_multiplicator => "1111011100110001",
            data_re_out => mul_re_out(963),
            data_im_out => mul_im_out(963)
        );

 
    UMUL_964 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(964),
            data_im_in => first_stage_im_out(964),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(964),
            data_im_out => mul_im_out(964)
        );

 
    UMUL_965 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(965),
            data_im_in => first_stage_im_out(965),
            re_multiplicator => "0011111001010000", --- 0.9736328125 + j-0.228088378906
            im_multiplicator => "1111000101100111",
            data_re_out => mul_re_out(965),
            data_im_out => mul_im_out(965)
        );

 
    UMUL_966 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(966),
            data_im_in => first_stage_im_out(966),
            re_multiplicator => "0011110110010011", --- 0.962097167969 + j-0.272644042969
            im_multiplicator => "1110111010001101",
            data_re_out => mul_re_out(966),
            data_im_out => mul_im_out(966)
        );

 
    UMUL_967 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(967),
            data_im_in => first_stage_im_out(967),
            re_multiplicator => "0011110010110101", --- 0.948547363281 + j-0.316589355469
            im_multiplicator => "1110101110111101",
            data_re_out => mul_re_out(967),
            data_im_out => mul_im_out(967)
        );

 
    UMUL_968 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(968),
            data_im_in => first_stage_im_out(968),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(968),
            data_im_out => mul_im_out(968)
        );

 
    UMUL_969 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(969),
            data_im_in => first_stage_im_out(969),
            re_multiplicator => "0011101010010111", --- 0.915466308594 + j-0.402404785156
            im_multiplicator => "1110011000111111",
            data_re_out => mul_re_out(969),
            data_im_out => mul_im_out(969)
        );

 
    UMUL_970 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(970),
            data_im_in => first_stage_im_out(970),
            re_multiplicator => "0011100101011000", --- 0.89599609375 + j-0.444091796875
            im_multiplicator => "1110001110010100",
            data_re_out => mul_re_out(970),
            data_im_out => mul_im_out(970)
        );

 
    UMUL_971 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(971),
            data_im_in => first_stage_im_out(971),
            re_multiplicator => "0011011111111001", --- 0.874572753906 + j-0.48486328125
            im_multiplicator => "1110000011111000",
            data_re_out => mul_re_out(971),
            data_im_out => mul_im_out(971)
        );

 
    UMUL_972 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(972),
            data_im_in => first_stage_im_out(972),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(972),
            data_im_out => mul_im_out(972)
        );

 
    UMUL_973 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(973),
            data_im_in => first_stage_im_out(973),
            re_multiplicator => "0011010011100010", --- 0.826293945312 + j-0.563171386719
            im_multiplicator => "1101101111110101",
            data_re_out => mul_re_out(973),
            data_im_out => mul_im_out(973)
        );

 
    UMUL_974 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(974),
            data_im_in => first_stage_im_out(974),
            re_multiplicator => "0011001100101100", --- 0.799560546875 + j-0.600646972656
            im_multiplicator => "1101100110001111",
            data_re_out => mul_re_out(974),
            data_im_out => mul_im_out(974)
        );

 
    UMUL_975 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(975),
            data_im_in => first_stage_im_out(975),
            re_multiplicator => "0011000101011001", --- 0.771057128906 + j-0.636779785156
            im_multiplicator => "1101011100111111",
            data_re_out => mul_re_out(975),
            data_im_out => mul_im_out(975)
        );

 
    UMUL_976 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(976),
            data_im_in => first_stage_im_out(976),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(976),
            data_im_out => mul_im_out(976)
        );

 
    UMUL_977 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(977),
            data_im_in => first_stage_im_out(977),
            re_multiplicator => "0010110101100101", --- 0.709289550781 + j-0.704956054688
            im_multiplicator => "1101001011100010",
            data_re_out => mul_re_out(977),
            data_im_out => mul_im_out(977)
        );

 
    UMUL_978 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(978),
            data_im_in => first_stage_im_out(978),
            re_multiplicator => "0010101101000101", --- 0.676086425781 + j-0.73681640625
            im_multiplicator => "1101000011011000",
            data_re_out => mul_re_out(978),
            data_im_out => mul_im_out(978)
        );

 
    UMUL_979 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(979),
            data_im_in => first_stage_im_out(979),
            re_multiplicator => "0010100100001110", --- 0.641479492188 + j-0.767150878906
            im_multiplicator => "1100111011100111",
            data_re_out => mul_re_out(979),
            data_im_out => mul_im_out(979)
        );

 
    UMUL_980 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(980),
            data_im_in => first_stage_im_out(980),
            re_multiplicator => "0010011011000001", --- 0.605529785156 + j-0.795837402344
            im_multiplicator => "1100110100010001",
            data_re_out => mul_re_out(980),
            data_im_out => mul_im_out(980)
        );

 
    UMUL_981 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(981),
            data_im_in => first_stage_im_out(981),
            re_multiplicator => "0010010001011110", --- 0.568237304688 + j-0.822875976562
            im_multiplicator => "1100101101010110",
            data_re_out => mul_re_out(981),
            data_im_out => mul_im_out(981)
        );

 
    UMUL_982 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(982),
            data_im_in => first_stage_im_out(982),
            re_multiplicator => "0010000111101000", --- 0.52978515625 + j-0.84814453125
            im_multiplicator => "1100100110111000",
            data_re_out => mul_re_out(982),
            data_im_out => mul_im_out(982)
        );

 
    UMUL_983 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(983),
            data_im_in => first_stage_im_out(983),
            re_multiplicator => "0001111101100000", --- 0.490234375 + j-0.87158203125
            im_multiplicator => "1100100000111000",
            data_re_out => mul_re_out(983),
            data_im_out => mul_im_out(983)
        );

 
    UMUL_984 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(984),
            data_im_in => first_stage_im_out(984),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(984),
            data_im_out => mul_im_out(984)
        );

 
    UMUL_985 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(985),
            data_im_in => first_stage_im_out(985),
            re_multiplicator => "0001101000011101", --- 0.408020019531 + j-0.912963867188
            im_multiplicator => "1100010110010010",
            data_re_out => mul_re_out(985),
            data_im_out => mul_im_out(985)
        );

 
    UMUL_986 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(986),
            data_im_in => first_stage_im_out(986),
            re_multiplicator => "0001011101100110", --- 0.365600585938 + j-0.930786132812
            im_multiplicator => "1100010001101110",
            data_re_out => mul_re_out(986),
            data_im_out => mul_im_out(986)
        );

 
    UMUL_987 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(987),
            data_im_in => first_stage_im_out(987),
            re_multiplicator => "0001010010100010", --- 0.322387695312 + j-0.946594238281
            im_multiplicator => "1100001101101011",
            data_re_out => mul_re_out(987),
            data_im_out => mul_im_out(987)
        );

 
    UMUL_988 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(988),
            data_im_in => first_stage_im_out(988),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(988),
            data_im_out => mul_im_out(988)
        );

 
    UMUL_989 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(989),
            data_im_in => first_stage_im_out(989),
            re_multiplicator => "0000111011111011", --- 0.234069824219 + j-0.972229003906
            im_multiplicator => "1100000111000111",
            data_re_out => mul_re_out(989),
            data_im_out => mul_im_out(989)
        );

 
    UMUL_990 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(990),
            data_im_in => first_stage_im_out(990),
            re_multiplicator => "0000110000011010", --- 0.189086914062 + j-0.98193359375
            im_multiplicator => "1100000100101000",
            data_re_out => mul_re_out(990),
            data_im_out => mul_im_out(990)
        );

 
    UMUL_991 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(991),
            data_im_in => first_stage_im_out(991),
            re_multiplicator => "0000100100110010", --- 0.143676757812 + j-0.989624023438
            im_multiplicator => "1100000010101010",
            data_re_out => mul_re_out(991),
            data_im_out => mul_im_out(991)
        );

 
    UMUL_992 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(992),
            data_im_in => first_stage_im_out(992),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(992),
            data_im_out => mul_im_out(992)
        );

 
    UMUL_993 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(993),
            data_im_in => first_stage_im_out(993),
            re_multiplicator => "0000001101010110", --- 0.0521240234375 + j-0.998657226562
            im_multiplicator => "1100000000010110",
            data_re_out => mul_re_out(993),
            data_im_out => mul_im_out(993)
        );

 
    UMUL_994 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(994),
            data_im_in => first_stage_im_out(994),
            re_multiplicator => "0000000001100101", --- 0.00616455078125 + j-1.0
            im_multiplicator => "1100000000000000",
            data_re_out => mul_re_out(994),
            data_im_out => mul_im_out(994)
        );

 
    UMUL_995 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(995),
            data_im_in => first_stage_im_out(995),
            re_multiplicator => "1111110101110011", --- -0.0398559570312 + j-0.999206542969
            im_multiplicator => "1100000000001101",
            data_re_out => mul_re_out(995),
            data_im_out => mul_im_out(995)
        );

 
    UMUL_996 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(996),
            data_im_in => first_stage_im_out(996),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(996),
            data_im_out => mul_im_out(996)
        );

 
    UMUL_997 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(997),
            data_im_in => first_stage_im_out(997),
            re_multiplicator => "1111011110010101", --- -0.131530761719 + j-0.991333007812
            im_multiplicator => "1100000010001110",
            data_re_out => mul_re_out(997),
            data_im_out => mul_im_out(997)
        );

 
    UMUL_998 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(998),
            data_im_in => first_stage_im_out(998),
            re_multiplicator => "1111010010101100", --- -0.177001953125 + j-0.984191894531
            im_multiplicator => "1100000100000011",
            data_re_out => mul_re_out(998),
            data_im_out => mul_im_out(998)
        );

 
    UMUL_999 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(999),
            data_im_in => first_stage_im_out(999),
            re_multiplicator => "1111000111001001", --- -0.222106933594 + j-0.975036621094
            im_multiplicator => "1100000110011001",
            data_re_out => mul_re_out(999),
            data_im_out => mul_im_out(999)
        );

 
    UMUL_1000 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1000),
            data_im_in => first_stage_im_out(1000),
            re_multiplicator => "1110111011101110", --- -0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(1000),
            data_im_out => mul_im_out(1000)
        );

 
    UMUL_1001 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1001),
            data_im_in => first_stage_im_out(1001),
            re_multiplicator => "1110110000011100", --- -0.310791015625 + j-0.950500488281
            im_multiplicator => "1100001100101011",
            data_re_out => mul_re_out(1001),
            data_im_out => mul_im_out(1001)
        );

 
    UMUL_1002 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1002),
            data_im_in => first_stage_im_out(1002),
            re_multiplicator => "1110100101010101", --- -0.354187011719 + j-0.935180664062
            im_multiplicator => "1100010000100110",
            data_re_out => mul_re_out(1002),
            data_im_out => mul_im_out(1002)
        );

 
    UMUL_1003 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1003),
            data_im_in => first_stage_im_out(1003),
            re_multiplicator => "1110011010011011", --- -0.396789550781 + j-0.917907714844
            im_multiplicator => "1100010101000001",
            data_re_out => mul_re_out(1003),
            data_im_out => mul_im_out(1003)
        );

 
    UMUL_1004 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1004),
            data_im_in => first_stage_im_out(1004),
            re_multiplicator => "1110001111101110", --- -0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(1004),
            data_im_out => mul_im_out(1004)
        );

 
    UMUL_1005 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1005),
            data_im_in => first_stage_im_out(1005),
            re_multiplicator => "1110000101010000", --- -0.4794921875 + j-0.877563476562
            im_multiplicator => "1100011111010110",
            data_re_out => mul_re_out(1005),
            data_im_out => mul_im_out(1005)
        );

 
    UMUL_1006 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1006),
            data_im_in => first_stage_im_out(1006),
            re_multiplicator => "1101111011000011", --- -0.519348144531 + j-0.854553222656
            im_multiplicator => "1100100101001111",
            data_re_out => mul_re_out(1006),
            data_im_out => mul_im_out(1006)
        );

 
    UMUL_1007 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1007),
            data_im_in => first_stage_im_out(1007),
            re_multiplicator => "1101110001001000", --- -0.55810546875 + j-0.829772949219
            im_multiplicator => "1100101011100101",
            data_re_out => mul_re_out(1007),
            data_im_out => mul_im_out(1007)
        );

 
    UMUL_1008 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1008),
            data_im_in => first_stage_im_out(1008),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(1008),
            data_im_out => mul_im_out(1008)
        );

 
    UMUL_1009 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1009),
            data_im_in => first_stage_im_out(1009),
            re_multiplicator => "1101011110001101", --- -0.632019042969 + j-0.774963378906
            im_multiplicator => "1100111001100111",
            data_re_out => mul_re_out(1009),
            data_im_out => mul_im_out(1009)
        );

 
    UMUL_1010 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1010),
            data_im_in => first_stage_im_out(1010),
            re_multiplicator => "1101010101010000", --- -0.6669921875 + j-0.745056152344
            im_multiplicator => "1101000001010001",
            data_re_out => mul_re_out(1010),
            data_im_out => mul_im_out(1010)
        );

 
    UMUL_1011 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1011),
            data_im_in => first_stage_im_out(1011),
            re_multiplicator => "1101001100101010", --- -0.700561523438 + j-0.713562011719
            im_multiplicator => "1101001001010101",
            data_re_out => mul_re_out(1011),
            data_im_out => mul_im_out(1011)
        );

 
    UMUL_1012 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1012),
            data_im_in => first_stage_im_out(1012),
            re_multiplicator => "1101000100011100", --- -0.732666015625 + j-0.680603027344
            im_multiplicator => "1101010001110001",
            data_re_out => mul_re_out(1012),
            data_im_out => mul_im_out(1012)
        );

 
    UMUL_1013 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1013),
            data_im_in => first_stage_im_out(1013),
            re_multiplicator => "1100111100101000", --- -0.76318359375 + j-0.646179199219
            im_multiplicator => "1101011010100101",
            data_re_out => mul_re_out(1013),
            data_im_out => mul_im_out(1013)
        );

 
    UMUL_1014 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1014),
            data_im_in => first_stage_im_out(1014),
            re_multiplicator => "1100110101001110", --- -0.792114257812 + j-0.610412597656
            im_multiplicator => "1101100011101111",
            data_re_out => mul_re_out(1014),
            data_im_out => mul_im_out(1014)
        );

 
    UMUL_1015 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1015),
            data_im_in => first_stage_im_out(1015),
            re_multiplicator => "1100101110010000", --- -0.8193359375 + j-0.573303222656
            im_multiplicator => "1101101101001111",
            data_re_out => mul_re_out(1015),
            data_im_out => mul_im_out(1015)
        );

 
    UMUL_1016 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1016),
            data_im_in => first_stage_im_out(1016),
            re_multiplicator => "1100100111101110", --- -0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(1016),
            data_im_out => mul_im_out(1016)
        );

 
    UMUL_1017 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1017),
            data_im_in => first_stage_im_out(1017),
            re_multiplicator => "1100100001101001", --- -0.868591308594 + j-0.495544433594
            im_multiplicator => "1110000001001001",
            data_re_out => mul_re_out(1017),
            data_im_out => mul_im_out(1017)
        );

 
    UMUL_1018 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1018),
            data_im_in => first_stage_im_out(1018),
            re_multiplicator => "1100011100000011", --- -0.890441894531 + j-0.455078125
            im_multiplicator => "1110001011100000",
            data_re_out => mul_re_out(1018),
            data_im_out => mul_im_out(1018)
        );

 
    UMUL_1019 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1019),
            data_im_in => first_stage_im_out(1019),
            re_multiplicator => "1100010110111011", --- -0.910461425781 + j-0.413635253906
            im_multiplicator => "1110010110000111",
            data_re_out => mul_re_out(1019),
            data_im_out => mul_im_out(1019)
        );

 
    UMUL_1020 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1020),
            data_im_in => first_stage_im_out(1020),
            re_multiplicator => "1100010010010011", --- -0.928527832031 + j-0.371337890625
            im_multiplicator => "1110100000111100",
            data_re_out => mul_re_out(1020),
            data_im_out => mul_im_out(1020)
        );

 
    UMUL_1021 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1021),
            data_im_in => first_stage_im_out(1021),
            re_multiplicator => "1100001110001100", --- -0.944580078125 + j-0.328186035156
            im_multiplicator => "1110101011111111",
            data_re_out => mul_re_out(1021),
            data_im_out => mul_im_out(1021)
        );

 
    UMUL_1022 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1022),
            data_im_in => first_stage_im_out(1022),
            re_multiplicator => "1100001010100101", --- -0.958679199219 + j-0.284423828125
            im_multiplicator => "1110110111001100",
            data_re_out => mul_re_out(1022),
            data_im_out => mul_im_out(1022)
        );

 
    UMUL_1023 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1023),
            data_im_in => first_stage_im_out(1023),
            re_multiplicator => "1100000111011111", --- -0.970764160156 + j-0.239990234375
            im_multiplicator => "1111000010100100",
            data_re_out => mul_re_out(1023),
            data_im_out => mul_im_out(1023)
        );

 
    UMUL_1024 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1024),
            data_im_in => first_stage_im_out(1024),
            data_re_out => mul_re_out(1024),
            data_im_out => mul_im_out(1024)
        );

 
    UMUL_1025 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1025),
            data_im_in => first_stage_im_out(1025),
            re_multiplicator => "0011111111101100", --- 0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(1025),
            data_im_out => mul_im_out(1025)
        );

 
    UMUL_1026 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1026),
            data_im_in => first_stage_im_out(1026),
            re_multiplicator => "0011111110110001", --- 0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(1026),
            data_im_out => mul_im_out(1026)
        );

 
    UMUL_1027 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1027),
            data_im_in => first_stage_im_out(1027),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(1027),
            data_im_out => mul_im_out(1027)
        );

 
    UMUL_1028 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1028),
            data_im_in => first_stage_im_out(1028),
            re_multiplicator => "0011111011000101", --- 0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(1028),
            data_im_out => mul_im_out(1028)
        );

 
    UMUL_1029 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1029),
            data_im_in => first_stage_im_out(1029),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(1029),
            data_im_out => mul_im_out(1029)
        );

 
    UMUL_1030 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1030),
            data_im_in => first_stage_im_out(1030),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(1030),
            data_im_out => mul_im_out(1030)
        );

 
    UMUL_1031 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1031),
            data_im_in => first_stage_im_out(1031),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(1031),
            data_im_out => mul_im_out(1031)
        );

 
    UMUL_1032 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1032),
            data_im_in => first_stage_im_out(1032),
            re_multiplicator => "0011101100100001", --- 0.923889160156 + j-0.382690429688
            im_multiplicator => "1110011110000010",
            data_re_out => mul_re_out(1032),
            data_im_out => mul_im_out(1032)
        );

 
    UMUL_1033 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1033),
            data_im_in => first_stage_im_out(1033),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(1033),
            data_im_out => mul_im_out(1033)
        );

 
    UMUL_1034 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1034),
            data_im_in => first_stage_im_out(1034),
            re_multiplicator => "0011100001110001", --- 0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(1034),
            data_im_out => mul_im_out(1034)
        );

 
    UMUL_1035 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1035),
            data_im_in => first_stage_im_out(1035),
            re_multiplicator => "0011011011100101", --- 0.857727050781 + j-0.514099121094
            im_multiplicator => "1101111100011001",
            data_re_out => mul_re_out(1035),
            data_im_out => mul_im_out(1035)
        );

 
    UMUL_1036 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1036),
            data_im_in => first_stage_im_out(1036),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(1036),
            data_im_out => mul_im_out(1036)
        );

 
    UMUL_1037 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1037),
            data_im_in => first_stage_im_out(1037),
            re_multiplicator => "0011001101101000", --- 0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(1037),
            data_im_out => mul_im_out(1037)
        );

 
    UMUL_1038 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1038),
            data_im_in => first_stage_im_out(1038),
            re_multiplicator => "0011000101111001", --- 0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(1038),
            data_im_out => mul_im_out(1038)
        );

 
    UMUL_1039 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1039),
            data_im_in => first_stage_im_out(1039),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(1039),
            data_im_out => mul_im_out(1039)
        );

 
    UMUL_1040 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1040),
            data_im_in => first_stage_im_out(1040),
            re_multiplicator => "0010110101000001", --- 0.707092285156 + j-0.707092285156
            im_multiplicator => "1101001010111111",
            data_re_out => mul_re_out(1040),
            data_im_out => mul_im_out(1040)
        );

 
    UMUL_1041 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1041),
            data_im_in => first_stage_im_out(1041),
            re_multiplicator => "0010101011111011", --- 0.671569824219 + j-0.740966796875
            im_multiplicator => "1101000010010100",
            data_re_out => mul_re_out(1041),
            data_im_out => mul_im_out(1041)
        );

 
    UMUL_1042 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1042),
            data_im_in => first_stage_im_out(1042),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(1042),
            data_im_out => mul_im_out(1042)
        );

 
    UMUL_1043 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1043),
            data_im_in => first_stage_im_out(1043),
            re_multiplicator => "0010011000100000", --- 0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(1043),
            data_im_out => mul_im_out(1043)
        );

 
    UMUL_1044 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1044),
            data_im_in => first_stage_im_out(1044),
            re_multiplicator => "0010001110001110", --- 0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(1044),
            data_im_out => mul_im_out(1044)
        );

 
    UMUL_1045 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1045),
            data_im_in => first_stage_im_out(1045),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(1045),
            data_im_out => mul_im_out(1045)
        );

 
    UMUL_1046 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1046),
            data_im_in => first_stage_im_out(1046),
            re_multiplicator => "0001111000101011", --- 0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(1046),
            data_im_out => mul_im_out(1046)
        );

 
    UMUL_1047 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1047),
            data_im_in => first_stage_im_out(1047),
            re_multiplicator => "0001101101011101", --- 0.427551269531 + j-0.903991699219
            im_multiplicator => "1100011000100101",
            data_re_out => mul_re_out(1047),
            data_im_out => mul_im_out(1047)
        );

 
    UMUL_1048 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1048),
            data_im_in => first_stage_im_out(1048),
            re_multiplicator => "0001100001111110", --- 0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(1048),
            data_im_out => mul_im_out(1048)
        );

 
    UMUL_1049 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1049),
            data_im_in => first_stage_im_out(1049),
            re_multiplicator => "0001010110010000", --- 0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(1049),
            data_im_out => mul_im_out(1049)
        );

 
    UMUL_1050 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1050),
            data_im_in => first_stage_im_out(1050),
            re_multiplicator => "0001001010010100", --- 0.290283203125 + j-0.956970214844
            im_multiplicator => "1100001011000001",
            data_re_out => mul_re_out(1050),
            data_im_out => mul_im_out(1050)
        );

 
    UMUL_1051 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1051),
            data_im_in => first_stage_im_out(1051),
            re_multiplicator => "0000111110001101", --- 0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(1051),
            data_im_out => mul_im_out(1051)
        );

 
    UMUL_1052 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1052),
            data_im_in => first_stage_im_out(1052),
            re_multiplicator => "0000110001111100", --- 0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(1052),
            data_im_out => mul_im_out(1052)
        );

 
    UMUL_1053 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1053),
            data_im_in => first_stage_im_out(1053),
            re_multiplicator => "0000100101100100", --- 0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(1053),
            data_im_out => mul_im_out(1053)
        );

 
    UMUL_1054 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1054),
            data_im_in => first_stage_im_out(1054),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(1054),
            data_im_out => mul_im_out(1054)
        );

 
    UMUL_1055 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1055),
            data_im_in => first_stage_im_out(1055),
            re_multiplicator => "0000001100100100", --- 0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(1055),
            data_im_out => mul_im_out(1055)
        );

 
    UMUL_1056 : multiplier_mulminusj
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1056),
            data_im_in => first_stage_im_out(1056),
            data_re_out => mul_re_out(1056),
            data_im_out => mul_im_out(1056)
        );

 
    UMUL_1057 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1057),
            data_im_in => first_stage_im_out(1057),
            re_multiplicator => "1111110011011100", --- -0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(1057),
            data_im_out => mul_im_out(1057)
        );

 
    UMUL_1058 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1058),
            data_im_in => first_stage_im_out(1058),
            re_multiplicator => "1111100110111010", --- -0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(1058),
            data_im_out => mul_im_out(1058)
        );

 
    UMUL_1059 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1059),
            data_im_in => first_stage_im_out(1059),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(1059),
            data_im_out => mul_im_out(1059)
        );

 
    UMUL_1060 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1060),
            data_im_in => first_stage_im_out(1060),
            re_multiplicator => "1111001110000100", --- -0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(1060),
            data_im_out => mul_im_out(1060)
        );

 
    UMUL_1061 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1061),
            data_im_in => first_stage_im_out(1061),
            re_multiplicator => "1111000001110011", --- -0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(1061),
            data_im_out => mul_im_out(1061)
        );

 
    UMUL_1062 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1062),
            data_im_in => first_stage_im_out(1062),
            re_multiplicator => "1110110101101100", --- -0.290283203125 + j-0.956970214844
            im_multiplicator => "1100001011000001",
            data_re_out => mul_re_out(1062),
            data_im_out => mul_im_out(1062)
        );

 
    UMUL_1063 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1063),
            data_im_in => first_stage_im_out(1063),
            re_multiplicator => "1110101001110000", --- -0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(1063),
            data_im_out => mul_im_out(1063)
        );

 
    UMUL_1064 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1064),
            data_im_in => first_stage_im_out(1064),
            re_multiplicator => "1110011110000010", --- -0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(1064),
            data_im_out => mul_im_out(1064)
        );

 
    UMUL_1065 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1065),
            data_im_in => first_stage_im_out(1065),
            re_multiplicator => "1110010010100011", --- -0.427551269531 + j-0.903991699219
            im_multiplicator => "1100011000100101",
            data_re_out => mul_re_out(1065),
            data_im_out => mul_im_out(1065)
        );

 
    UMUL_1066 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1066),
            data_im_in => first_stage_im_out(1066),
            re_multiplicator => "1110000111010101", --- -0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(1066),
            data_im_out => mul_im_out(1066)
        );

 
    UMUL_1067 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1067),
            data_im_in => first_stage_im_out(1067),
            re_multiplicator => "1101111100011001", --- -0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(1067),
            data_im_out => mul_im_out(1067)
        );

 
    UMUL_1068 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1068),
            data_im_in => first_stage_im_out(1068),
            re_multiplicator => "1101110001110010", --- -0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(1068),
            data_im_out => mul_im_out(1068)
        );

 
    UMUL_1069 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1069),
            data_im_in => first_stage_im_out(1069),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(1069),
            data_im_out => mul_im_out(1069)
        );

 
    UMUL_1070 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1070),
            data_im_in => first_stage_im_out(1070),
            re_multiplicator => "1101011101100110", --- -0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(1070),
            data_im_out => mul_im_out(1070)
        );

 
    UMUL_1071 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1071),
            data_im_in => first_stage_im_out(1071),
            re_multiplicator => "1101010100000101", --- -0.671569824219 + j-0.740966796875
            im_multiplicator => "1101000010010100",
            data_re_out => mul_re_out(1071),
            data_im_out => mul_im_out(1071)
        );

 
    UMUL_1072 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1072),
            data_im_in => first_stage_im_out(1072),
            re_multiplicator => "1101001010111111", --- -0.707092285156 + j-0.707092285156
            im_multiplicator => "1101001010111111",
            data_re_out => mul_re_out(1072),
            data_im_out => mul_im_out(1072)
        );

 
    UMUL_1073 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1073),
            data_im_in => first_stage_im_out(1073),
            re_multiplicator => "1101000010010100", --- -0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(1073),
            data_im_out => mul_im_out(1073)
        );

 
    UMUL_1074 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1074),
            data_im_in => first_stage_im_out(1074),
            re_multiplicator => "1100111010000111", --- -0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(1074),
            data_im_out => mul_im_out(1074)
        );

 
    UMUL_1075 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1075),
            data_im_in => first_stage_im_out(1075),
            re_multiplicator => "1100110010011000", --- -0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(1075),
            data_im_out => mul_im_out(1075)
        );

 
    UMUL_1076 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1076),
            data_im_in => first_stage_im_out(1076),
            re_multiplicator => "1100101011001001", --- -0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(1076),
            data_im_out => mul_im_out(1076)
        );

 
    UMUL_1077 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1077),
            data_im_in => first_stage_im_out(1077),
            re_multiplicator => "1100100100011011", --- -0.857727050781 + j-0.514099121094
            im_multiplicator => "1101111100011001",
            data_re_out => mul_re_out(1077),
            data_im_out => mul_im_out(1077)
        );

 
    UMUL_1078 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1078),
            data_im_in => first_stage_im_out(1078),
            re_multiplicator => "1100011110001111", --- -0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(1078),
            data_im_out => mul_im_out(1078)
        );

 
    UMUL_1079 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1079),
            data_im_in => first_stage_im_out(1079),
            re_multiplicator => "1100011000100101", --- -0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(1079),
            data_im_out => mul_im_out(1079)
        );

 
    UMUL_1080 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1080),
            data_im_in => first_stage_im_out(1080),
            re_multiplicator => "1100010011011111", --- -0.923889160156 + j-0.382690429688
            im_multiplicator => "1110011110000010",
            data_re_out => mul_re_out(1080),
            data_im_out => mul_im_out(1080)
        );

 
    UMUL_1081 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1081),
            data_im_in => first_stage_im_out(1081),
            re_multiplicator => "1100001110111110", --- -0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(1081),
            data_im_out => mul_im_out(1081)
        );

 
    UMUL_1082 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1082),
            data_im_in => first_stage_im_out(1082),
            re_multiplicator => "1100001011000001", --- -0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(1082),
            data_im_out => mul_im_out(1082)
        );

 
    UMUL_1083 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1083),
            data_im_in => first_stage_im_out(1083),
            re_multiplicator => "1100000111101011", --- -0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(1083),
            data_im_out => mul_im_out(1083)
        );

 
    UMUL_1084 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1084),
            data_im_in => first_stage_im_out(1084),
            re_multiplicator => "1100000100111011", --- -0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(1084),
            data_im_out => mul_im_out(1084)
        );

 
    UMUL_1085 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1085),
            data_im_in => first_stage_im_out(1085),
            re_multiplicator => "1100000010110001", --- -0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(1085),
            data_im_out => mul_im_out(1085)
        );

 
    UMUL_1086 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1086),
            data_im_in => first_stage_im_out(1086),
            re_multiplicator => "1100000001001111", --- -0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(1086),
            data_im_out => mul_im_out(1086)
        );

 
    UMUL_1087 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1087),
            data_im_in => first_stage_im_out(1087),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(1087),
            data_im_out => mul_im_out(1087)
        );

 
    UMUL_1088 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1088),
            data_im_in => first_stage_im_out(1088),
            data_re_out => mul_re_out(1088),
            data_im_out => mul_im_out(1088)
        );

 
    UMUL_1089 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1089),
            data_im_in => first_stage_im_out(1089),
            re_multiplicator => "0011111111101010", --- 0.998657226562 + j-0.0521240234375
            im_multiplicator => "1111110010101010",
            data_re_out => mul_re_out(1089),
            data_im_out => mul_im_out(1089)
        );

 
    UMUL_1090 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1090),
            data_im_in => first_stage_im_out(1090),
            re_multiplicator => "0011111110100111", --- 0.994567871094 + j-0.104125976562
            im_multiplicator => "1111100101010110",
            data_re_out => mul_re_out(1090),
            data_im_out => mul_im_out(1090)
        );

 
    UMUL_1091 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1091),
            data_im_in => first_stage_im_out(1091),
            re_multiplicator => "0011111100111000", --- 0.98779296875 + j-0.155822753906
            im_multiplicator => "1111011000000111",
            data_re_out => mul_re_out(1091),
            data_im_out => mul_im_out(1091)
        );

 
    UMUL_1092 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1092),
            data_im_in => first_stage_im_out(1092),
            re_multiplicator => "0011111010011101", --- 0.978332519531 + j-0.207092285156
            im_multiplicator => "1111001010111111",
            data_re_out => mul_re_out(1092),
            data_im_out => mul_im_out(1092)
        );

 
    UMUL_1093 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1093),
            data_im_in => first_stage_im_out(1093),
            re_multiplicator => "0011110111010110", --- 0.966186523438 + j-0.2578125
            im_multiplicator => "1110111110000000",
            data_re_out => mul_re_out(1093),
            data_im_out => mul_im_out(1093)
        );

 
    UMUL_1094 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1094),
            data_im_in => first_stage_im_out(1094),
            re_multiplicator => "0011110011100100", --- 0.951416015625 + j-0.307861328125
            im_multiplicator => "1110110001001100",
            data_re_out => mul_re_out(1094),
            data_im_out => mul_im_out(1094)
        );

 
    UMUL_1095 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1095),
            data_im_in => first_stage_im_out(1095),
            re_multiplicator => "0011101111001000", --- 0.93408203125 + j-0.357055664062
            im_multiplicator => "1110100100100110",
            data_re_out => mul_re_out(1095),
            data_im_out => mul_im_out(1095)
        );

 
    UMUL_1096 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1096),
            data_im_in => first_stage_im_out(1096),
            re_multiplicator => "0011101010000010", --- 0.914184570312 + j-0.405212402344
            im_multiplicator => "1110011000010001",
            data_re_out => mul_re_out(1096),
            data_im_out => mul_im_out(1096)
        );

 
    UMUL_1097 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1097),
            data_im_in => first_stage_im_out(1097),
            re_multiplicator => "0011100100010100", --- 0.891845703125 + j-0.452331542969
            im_multiplicator => "1110001100001101",
            data_re_out => mul_re_out(1097),
            data_im_out => mul_im_out(1097)
        );

 
    UMUL_1098 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1098),
            data_im_in => first_stage_im_out(1098),
            re_multiplicator => "0011011101111110", --- 0.867065429688 + j-0.498229980469
            im_multiplicator => "1110000000011101",
            data_re_out => mul_re_out(1098),
            data_im_out => mul_im_out(1098)
        );

 
    UMUL_1099 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1099),
            data_im_in => first_stage_im_out(1099),
            re_multiplicator => "0011010111000001", --- 0.839904785156 + j-0.542724609375
            im_multiplicator => "1101110101000100",
            data_re_out => mul_re_out(1099),
            data_im_out => mul_im_out(1099)
        );

 
    UMUL_1100 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1100),
            data_im_in => first_stage_im_out(1100),
            re_multiplicator => "0011001111011111", --- 0.810485839844 + j-0.585815429688
            im_multiplicator => "1101101010000010",
            data_re_out => mul_re_out(1100),
            data_im_out => mul_im_out(1100)
        );

 
    UMUL_1101 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1101),
            data_im_in => first_stage_im_out(1101),
            re_multiplicator => "0011000111011000", --- 0.77880859375 + j-0.627258300781
            im_multiplicator => "1101011111011011",
            data_re_out => mul_re_out(1101),
            data_im_out => mul_im_out(1101)
        );

 
    UMUL_1102 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1102),
            data_im_in => first_stage_im_out(1102),
            re_multiplicator => "0010111110101111", --- 0.745056152344 + j-0.6669921875
            im_multiplicator => "1101010101010000",
            data_re_out => mul_re_out(1102),
            data_im_out => mul_im_out(1102)
        );

 
    UMUL_1103 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1103),
            data_im_in => first_stage_im_out(1103),
            re_multiplicator => "0010110101100101", --- 0.709289550781 + j-0.704956054688
            im_multiplicator => "1101001011100010",
            data_re_out => mul_re_out(1103),
            data_im_out => mul_im_out(1103)
        );

 
    UMUL_1104 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1104),
            data_im_in => first_stage_im_out(1104),
            re_multiplicator => "0010101011111011", --- 0.671569824219 + j-0.740966796875
            im_multiplicator => "1101000010010100",
            data_re_out => mul_re_out(1104),
            data_im_out => mul_im_out(1104)
        );

 
    UMUL_1105 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1105),
            data_im_in => first_stage_im_out(1105),
            re_multiplicator => "0010100001110011", --- 0.632019042969 + j-0.774963378906
            im_multiplicator => "1100111001100111",
            data_re_out => mul_re_out(1105),
            data_im_out => mul_im_out(1105)
        );

 
    UMUL_1106 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1106),
            data_im_in => first_stage_im_out(1106),
            re_multiplicator => "0010010111001111", --- 0.590759277344 + j-0.806823730469
            im_multiplicator => "1100110001011101",
            data_re_out => mul_re_out(1106),
            data_im_out => mul_im_out(1106)
        );

 
    UMUL_1107 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1107),
            data_im_in => first_stage_im_out(1107),
            re_multiplicator => "0010001100010001", --- 0.547912597656 + j-0.836547851562
            im_multiplicator => "1100101001110110",
            data_re_out => mul_re_out(1107),
            data_im_out => mul_im_out(1107)
        );

 
    UMUL_1108 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1108),
            data_im_in => first_stage_im_out(1108),
            re_multiplicator => "0010000000111010", --- 0.503540039062 + j-0.863952636719
            im_multiplicator => "1100100010110101",
            data_re_out => mul_re_out(1108),
            data_im_out => mul_im_out(1108)
        );

 
    UMUL_1109 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1109),
            data_im_in => first_stage_im_out(1109),
            re_multiplicator => "0001110101001101", --- 0.457824707031 + j-0.889038085938
            im_multiplicator => "1100011100011010",
            data_re_out => mul_re_out(1109),
            data_im_out => mul_im_out(1109)
        );

 
    UMUL_1110 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1110),
            data_im_in => first_stage_im_out(1110),
            re_multiplicator => "0001101001001011", --- 0.410827636719 + j-0.911682128906
            im_multiplicator => "1100010110100111",
            data_re_out => mul_re_out(1110),
            data_im_out => mul_im_out(1110)
        );

 
    UMUL_1111 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1111),
            data_im_in => first_stage_im_out(1111),
            re_multiplicator => "0001011100110111", --- 0.362731933594 + j-0.931884765625
            im_multiplicator => "1100010001011100",
            data_re_out => mul_re_out(1111),
            data_im_out => mul_im_out(1111)
        );

 
    UMUL_1112 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1112),
            data_im_in => first_stage_im_out(1112),
            re_multiplicator => "0001010000010011", --- 0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(1112),
            data_im_out => mul_im_out(1112)
        );

 
    UMUL_1113 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1113),
            data_im_in => first_stage_im_out(1113),
            re_multiplicator => "0001000011100001", --- 0.263732910156 + j-0.964599609375
            im_multiplicator => "1100001001000100",
            data_re_out => mul_re_out(1113),
            data_im_out => mul_im_out(1113)
        );

 
    UMUL_1114 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1114),
            data_im_in => first_stage_im_out(1114),
            re_multiplicator => "0000110110100100", --- 0.213134765625 + j-0.97705078125
            im_multiplicator => "1100000101111000",
            data_re_out => mul_re_out(1114),
            data_im_out => mul_im_out(1114)
        );

 
    UMUL_1115 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1115),
            data_im_in => first_stage_im_out(1115),
            re_multiplicator => "0000101001011100", --- 0.161865234375 + j-0.98681640625
            im_multiplicator => "1100000011011000",
            data_re_out => mul_re_out(1115),
            data_im_out => mul_im_out(1115)
        );

 
    UMUL_1116 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1116),
            data_im_in => first_stage_im_out(1116),
            re_multiplicator => "0000011100001110", --- 0.110229492188 + j-0.993896484375
            im_multiplicator => "1100000001100100",
            data_re_out => mul_re_out(1116),
            data_im_out => mul_im_out(1116)
        );

 
    UMUL_1117 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1117),
            data_im_in => first_stage_im_out(1117),
            re_multiplicator => "0000001110111011", --- 0.0582885742188 + j-0.998291015625
            im_multiplicator => "1100000000011100",
            data_re_out => mul_re_out(1117),
            data_im_out => mul_im_out(1117)
        );

 
    UMUL_1118 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1118),
            data_im_in => first_stage_im_out(1118),
            re_multiplicator => "0000000001100101", --- 0.00616455078125 + j-1.0
            im_multiplicator => "1100000000000000",
            data_re_out => mul_re_out(1118),
            data_im_out => mul_im_out(1118)
        );

 
    UMUL_1119 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1119),
            data_im_in => first_stage_im_out(1119),
            re_multiplicator => "1111110100001110", --- -0.0460205078125 + j-0.998962402344
            im_multiplicator => "1100000000010001",
            data_re_out => mul_re_out(1119),
            data_im_out => mul_im_out(1119)
        );

 
    UMUL_1120 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1120),
            data_im_in => first_stage_im_out(1120),
            re_multiplicator => "1111100110111010", --- -0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(1120),
            data_im_out => mul_im_out(1120)
        );

 
    UMUL_1121 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1121),
            data_im_in => first_stage_im_out(1121),
            re_multiplicator => "1111011001101010", --- -0.149780273438 + j-0.988708496094
            im_multiplicator => "1100000010111001",
            data_re_out => mul_re_out(1121),
            data_im_out => mul_im_out(1121)
        );

 
    UMUL_1122 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1122),
            data_im_in => first_stage_im_out(1122),
            re_multiplicator => "1111001100100001", --- -0.201110839844 + j-0.979553222656
            im_multiplicator => "1100000101001111",
            data_re_out => mul_re_out(1122),
            data_im_out => mul_im_out(1122)
        );

 
    UMUL_1123 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1123),
            data_im_in => first_stage_im_out(1123),
            re_multiplicator => "1110111111100001", --- -0.251892089844 + j-0.9677734375
            im_multiplicator => "1100001000010000",
            data_re_out => mul_re_out(1123),
            data_im_out => mul_im_out(1123)
        );

 
    UMUL_1124 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1124),
            data_im_in => first_stage_im_out(1124),
            re_multiplicator => "1110110010101100", --- -0.302001953125 + j-0.953308105469
            im_multiplicator => "1100001011111101",
            data_re_out => mul_re_out(1124),
            data_im_out => mul_im_out(1124)
        );

 
    UMUL_1125 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1125),
            data_im_in => first_stage_im_out(1125),
            re_multiplicator => "1110100110000100", --- -0.351318359375 + j-0.936279296875
            im_multiplicator => "1100010000010100",
            data_re_out => mul_re_out(1125),
            data_im_out => mul_im_out(1125)
        );

 
    UMUL_1126 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1126),
            data_im_in => first_stage_im_out(1126),
            re_multiplicator => "1110011001101101", --- -0.399597167969 + j-0.916687011719
            im_multiplicator => "1100010101010101",
            data_re_out => mul_re_out(1126),
            data_im_out => mul_im_out(1126)
        );

 
    UMUL_1127 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1127),
            data_im_in => first_stage_im_out(1127),
            re_multiplicator => "1110001101100111", --- -0.446838378906 + j-0.894592285156
            im_multiplicator => "1100011010111111",
            data_re_out => mul_re_out(1127),
            data_im_out => mul_im_out(1127)
        );

 
    UMUL_1128 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1128),
            data_im_in => first_stage_im_out(1128),
            re_multiplicator => "1110000001110100", --- -0.492919921875 + j-0.8701171875
            im_multiplicator => "1100100001010000",
            data_re_out => mul_re_out(1128),
            data_im_out => mul_im_out(1128)
        );

 
    UMUL_1129 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1129),
            data_im_in => first_stage_im_out(1129),
            re_multiplicator => "1101110110011000", --- -0.53759765625 + j-0.843200683594
            im_multiplicator => "1100101000001001",
            data_re_out => mul_re_out(1129),
            data_im_out => mul_im_out(1129)
        );

 
    UMUL_1130 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1130),
            data_im_in => first_stage_im_out(1130),
            re_multiplicator => "1101101011010100", --- -0.580810546875 + j-0.814025878906
            im_multiplicator => "1100101111100111",
            data_re_out => mul_re_out(1130),
            data_im_out => mul_im_out(1130)
        );

 
    UMUL_1131 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1131),
            data_im_in => first_stage_im_out(1131),
            re_multiplicator => "1101100000101010", --- -0.622436523438 + j-0.782653808594
            im_multiplicator => "1100110111101001",
            data_re_out => mul_re_out(1131),
            data_im_out => mul_im_out(1131)
        );

 
    UMUL_1132 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1132),
            data_im_in => first_stage_im_out(1132),
            re_multiplicator => "1101010110011011", --- -0.662414550781 + j-0.749145507812
            im_multiplicator => "1101000000001110",
            data_re_out => mul_re_out(1132),
            data_im_out => mul_im_out(1132)
        );

 
    UMUL_1133 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1133),
            data_im_in => first_stage_im_out(1133),
            re_multiplicator => "1101001100101010", --- -0.700561523438 + j-0.713562011719
            im_multiplicator => "1101001001010101",
            data_re_out => mul_re_out(1133),
            data_im_out => mul_im_out(1133)
        );

 
    UMUL_1134 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1134),
            data_im_in => first_stage_im_out(1134),
            re_multiplicator => "1101000011011000", --- -0.73681640625 + j-0.676086425781
            im_multiplicator => "1101010010111011",
            data_re_out => mul_re_out(1134),
            data_im_out => mul_im_out(1134)
        );

 
    UMUL_1135 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1135),
            data_im_in => first_stage_im_out(1135),
            re_multiplicator => "1100111010100111", --- -0.771057128906 + j-0.636779785156
            im_multiplicator => "1101011100111111",
            data_re_out => mul_re_out(1135),
            data_im_out => mul_im_out(1135)
        );

 
    UMUL_1136 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1136),
            data_im_in => first_stage_im_out(1136),
            re_multiplicator => "1100110010011000", --- -0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(1136),
            data_im_out => mul_im_out(1136)
        );

 
    UMUL_1137 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1137),
            data_im_in => first_stage_im_out(1137),
            re_multiplicator => "1100101010101101", --- -0.833190917969 + j-0.553039550781
            im_multiplicator => "1101110010011011",
            data_re_out => mul_re_out(1137),
            data_im_out => mul_im_out(1137)
        );

 
    UMUL_1138 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1138),
            data_im_in => first_stage_im_out(1138),
            re_multiplicator => "1100100011101000", --- -0.86083984375 + j-0.508850097656
            im_multiplicator => "1101111101101111",
            data_re_out => mul_re_out(1138),
            data_im_out => mul_im_out(1138)
        );

 
    UMUL_1139 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1139),
            data_im_in => first_stage_im_out(1139),
            re_multiplicator => "1100011101001000", --- -0.88623046875 + j-0.463256835938
            im_multiplicator => "1110001001011010",
            data_re_out => mul_re_out(1139),
            data_im_out => mul_im_out(1139)
        );

 
    UMUL_1140 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1140),
            data_im_in => first_stage_im_out(1140),
            re_multiplicator => "1100010111010000", --- -0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(1140),
            data_im_out => mul_im_out(1140)
        );

 
    UMUL_1141 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1141),
            data_im_in => first_stage_im_out(1141),
            re_multiplicator => "1100010010000001", --- -0.929626464844 + j-0.368469238281
            im_multiplicator => "1110100001101011",
            data_re_out => mul_re_out(1141),
            data_im_out => mul_im_out(1141)
        );

 
    UMUL_1142 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1142),
            data_im_in => first_stage_im_out(1142),
            re_multiplicator => "1100001101011011", --- -0.947570800781 + j-0.319519042969
            im_multiplicator => "1110101110001101",
            data_re_out => mul_re_out(1142),
            data_im_out => mul_im_out(1142)
        );

 
    UMUL_1143 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1143),
            data_im_in => first_stage_im_out(1143),
            re_multiplicator => "1100001001011111", --- -0.962951660156 + j-0.269653320312
            im_multiplicator => "1110111010111110",
            data_re_out => mul_re_out(1143),
            data_im_out => mul_im_out(1143)
        );

 
    UMUL_1144 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1144),
            data_im_in => first_stage_im_out(1144),
            re_multiplicator => "1100000110001110", --- -0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(1144),
            data_im_out => mul_im_out(1144)
        );

 
    UMUL_1145 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1145),
            data_im_in => first_stage_im_out(1145),
            re_multiplicator => "1100000011101001", --- -0.985778808594 + j-0.16796875
            im_multiplicator => "1111010101000000",
            data_re_out => mul_re_out(1145),
            data_im_out => mul_im_out(1145)
        );

 
    UMUL_1146 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1146),
            data_im_in => first_stage_im_out(1146),
            re_multiplicator => "1100000001101111", --- -0.993225097656 + j-0.116333007812
            im_multiplicator => "1111100010001110",
            data_re_out => mul_re_out(1146),
            data_im_out => mul_im_out(1146)
        );

 
    UMUL_1147 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1147),
            data_im_in => first_stage_im_out(1147),
            re_multiplicator => "1100000000100010", --- -0.997924804688 + j-0.0643920898438
            im_multiplicator => "1111101111100001",
            data_re_out => mul_re_out(1147),
            data_im_out => mul_im_out(1147)
        );

 
    UMUL_1148 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1148),
            data_im_in => first_stage_im_out(1148),
            re_multiplicator => "1100000000000001", --- -0.999938964844 + j-0.0122680664062
            im_multiplicator => "1111111100110111",
            data_re_out => mul_re_out(1148),
            data_im_out => mul_im_out(1148)
        );

 
    UMUL_1149 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1149),
            data_im_in => first_stage_im_out(1149),
            re_multiplicator => "1100000000001101", --- -0.999206542969 + j0.0398559570312
            im_multiplicator => "0000001010001101",
            data_re_out => mul_re_out(1149),
            data_im_out => mul_im_out(1149)
        );

 
    UMUL_1150 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1150),
            data_im_in => first_stage_im_out(1150),
            re_multiplicator => "1100000001000101", --- -0.995788574219 + j0.0919189453125
            im_multiplicator => "0000010111100010",
            data_re_out => mul_re_out(1150),
            data_im_out => mul_im_out(1150)
        );

 
    UMUL_1151 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1151),
            data_im_in => first_stage_im_out(1151),
            re_multiplicator => "1100000010101010", --- -0.989624023438 + j0.143676757812
            im_multiplicator => "0000100100110010",
            data_re_out => mul_re_out(1151),
            data_im_out => mul_im_out(1151)
        );

 
    UMUL_1152 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1152),
            data_im_in => first_stage_im_out(1152),
            data_re_out => mul_re_out(1152),
            data_im_out => mul_im_out(1152)
        );

 
    UMUL_1153 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1153),
            data_im_in => first_stage_im_out(1153),
            re_multiplicator => "0011111111100111", --- 0.998474121094 + j-0.05517578125
            im_multiplicator => "1111110001111000",
            data_re_out => mul_re_out(1153),
            data_im_out => mul_im_out(1153)
        );

 
    UMUL_1154 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1154),
            data_im_in => first_stage_im_out(1154),
            re_multiplicator => "0011111110011100", --- 0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(1154),
            data_im_out => mul_im_out(1154)
        );

 
    UMUL_1155 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1155),
            data_im_in => first_stage_im_out(1155),
            re_multiplicator => "0011111100100000", --- 0.986328125 + j-0.164916992188
            im_multiplicator => "1111010101110010",
            data_re_out => mul_re_out(1155),
            data_im_out => mul_im_out(1155)
        );

 
    UMUL_1156 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1156),
            data_im_in => first_stage_im_out(1156),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(1156),
            data_im_out => mul_im_out(1156)
        );

 
    UMUL_1157 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1157),
            data_im_in => first_stage_im_out(1157),
            re_multiplicator => "0011110110010011", --- 0.962097167969 + j-0.272644042969
            im_multiplicator => "1110111010001101",
            data_re_out => mul_re_out(1157),
            data_im_out => mul_im_out(1157)
        );

 
    UMUL_1158 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1158),
            data_im_in => first_stage_im_out(1158),
            re_multiplicator => "0011110010000101", --- 0.945617675781 + j-0.325317382812
            im_multiplicator => "1110101100101110",
            data_re_out => mul_re_out(1158),
            data_im_out => mul_im_out(1158)
        );

 
    UMUL_1159 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1159),
            data_im_in => first_stage_im_out(1159),
            re_multiplicator => "0011101101000111", --- 0.926208496094 + j-0.377014160156
            im_multiplicator => "1110011111011111",
            data_re_out => mul_re_out(1159),
            data_im_out => mul_im_out(1159)
        );

 
    UMUL_1160 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1160),
            data_im_in => first_stage_im_out(1160),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(1160),
            data_im_out => mul_im_out(1160)
        );

 
    UMUL_1161 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1161),
            data_im_in => first_stage_im_out(1161),
            re_multiplicator => "0011100001000010", --- 0.879028320312 + j-0.476806640625
            im_multiplicator => "1110000101111100",
            data_re_out => mul_re_out(1161),
            data_im_out => mul_im_out(1161)
        );

 
    UMUL_1162 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1162),
            data_im_in => first_stage_im_out(1162),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(1162),
            data_im_out => mul_im_out(1162)
        );

 
    UMUL_1163 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1163),
            data_im_in => first_stage_im_out(1163),
            re_multiplicator => "0011010010001101", --- 0.821105957031 + j-0.57080078125
            im_multiplicator => "1101101101111000",
            data_re_out => mul_re_out(1163),
            data_im_out => mul_im_out(1163)
        );

 
    UMUL_1164 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1164),
            data_im_in => first_stage_im_out(1164),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(1164),
            data_im_out => mul_im_out(1164)
        );

 
    UMUL_1165 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1165),
            data_im_in => first_stage_im_out(1165),
            re_multiplicator => "0011000000110100", --- 0.753173828125 + j-0.657836914062
            im_multiplicator => "1101010111100110",
            data_re_out => mul_re_out(1165),
            data_im_out => mul_im_out(1165)
        );

 
    UMUL_1166 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1166),
            data_im_in => first_stage_im_out(1166),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(1166),
            data_im_out => mul_im_out(1166)
        );

 
    UMUL_1167 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1167),
            data_im_in => first_stage_im_out(1167),
            re_multiplicator => "0010101101000101", --- 0.676086425781 + j-0.73681640625
            im_multiplicator => "1101000011011000",
            data_re_out => mul_re_out(1167),
            data_im_out => mul_im_out(1167)
        );

 
    UMUL_1168 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1168),
            data_im_in => first_stage_im_out(1168),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(1168),
            data_im_out => mul_im_out(1168)
        );

 
    UMUL_1169 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1169),
            data_im_in => first_stage_im_out(1169),
            re_multiplicator => "0010010111001111", --- 0.590759277344 + j-0.806823730469
            im_multiplicator => "1100110001011101",
            data_re_out => mul_re_out(1169),
            data_im_out => mul_im_out(1169)
        );

 
    UMUL_1170 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1170),
            data_im_in => first_stage_im_out(1170),
            re_multiplicator => "0010001011100111", --- 0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(1170),
            data_im_out => mul_im_out(1170)
        );

 
    UMUL_1171 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1171),
            data_im_in => first_stage_im_out(1171),
            re_multiplicator => "0001111111100011", --- 0.498229980469 + j-0.867065429688
            im_multiplicator => "1100100010000010",
            data_re_out => mul_re_out(1171),
            data_im_out => mul_im_out(1171)
        );

 
    UMUL_1172 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1172),
            data_im_in => first_stage_im_out(1172),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(1172),
            data_im_out => mul_im_out(1172)
        );

 
    UMUL_1173 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1173),
            data_im_in => first_stage_im_out(1173),
            re_multiplicator => "0001100110010011", --- 0.399597167969 + j-0.916687011719
            im_multiplicator => "1100010101010101",
            data_re_out => mul_re_out(1173),
            data_im_out => mul_im_out(1173)
        );

 
    UMUL_1174 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1174),
            data_im_in => first_stage_im_out(1174),
            re_multiplicator => "0001011001001100", --- 0.348388671875 + j-0.937316894531
            im_multiplicator => "1100010000000011",
            data_re_out => mul_re_out(1174),
            data_im_out => mul_im_out(1174)
        );

 
    UMUL_1175 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1175),
            data_im_in => first_stage_im_out(1175),
            re_multiplicator => "0001001011110100", --- 0.296142578125 + j-0.955139160156
            im_multiplicator => "1100001011011111",
            data_re_out => mul_re_out(1175),
            data_im_out => mul_im_out(1175)
        );

 
    UMUL_1176 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1176),
            data_im_in => first_stage_im_out(1176),
            re_multiplicator => "0000111110001101", --- 0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(1176),
            data_im_out => mul_im_out(1176)
        );

 
    UMUL_1177 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1177),
            data_im_in => first_stage_im_out(1177),
            re_multiplicator => "0000110000011010", --- 0.189086914062 + j-0.98193359375
            im_multiplicator => "1100000100101000",
            data_re_out => mul_re_out(1177),
            data_im_out => mul_im_out(1177)
        );

 
    UMUL_1178 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1178),
            data_im_in => first_stage_im_out(1178),
            re_multiplicator => "0000100010011101", --- 0.134582519531 + j-0.990905761719
            im_multiplicator => "1100000010010101",
            data_re_out => mul_re_out(1178),
            data_im_out => mul_im_out(1178)
        );

 
    UMUL_1179 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1179),
            data_im_in => first_stage_im_out(1179),
            re_multiplicator => "0000010100011010", --- 0.0797119140625 + j-0.996826171875
            im_multiplicator => "1100000000110100",
            data_re_out => mul_re_out(1179),
            data_im_out => mul_im_out(1179)
        );

 
    UMUL_1180 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1180),
            data_im_in => first_stage_im_out(1180),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(1180),
            data_im_out => mul_im_out(1180)
        );

 
    UMUL_1181 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1181),
            data_im_in => first_stage_im_out(1181),
            re_multiplicator => "1111111000001001", --- -0.0307006835938 + j-0.99951171875
            im_multiplicator => "1100000000001000",
            data_re_out => mul_re_out(1181),
            data_im_out => mul_im_out(1181)
        );

 
    UMUL_1182 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1182),
            data_im_in => first_stage_im_out(1182),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(1182),
            data_im_out => mul_im_out(1182)
        );

 
    UMUL_1183 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1183),
            data_im_in => first_stage_im_out(1183),
            re_multiplicator => "1111011011111111", --- -0.140686035156 + j-0.990051269531
            im_multiplicator => "1100000010100011",
            data_re_out => mul_re_out(1183),
            data_im_out => mul_im_out(1183)
        );

 
    UMUL_1184 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1184),
            data_im_in => first_stage_im_out(1184),
            re_multiplicator => "1111001110000100", --- -0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(1184),
            data_im_out => mul_im_out(1184)
        );

 
    UMUL_1185 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1185),
            data_im_in => first_stage_im_out(1185),
            re_multiplicator => "1111000000010010", --- -0.248901367188 + j-0.968505859375
            im_multiplicator => "1100001000000100",
            data_re_out => mul_re_out(1185),
            data_im_out => mul_im_out(1185)
        );

 
    UMUL_1186 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1186),
            data_im_in => first_stage_im_out(1186),
            re_multiplicator => "1110110010101100", --- -0.302001953125 + j-0.953308105469
            im_multiplicator => "1100001011111101",
            data_re_out => mul_re_out(1186),
            data_im_out => mul_im_out(1186)
        );

 
    UMUL_1187 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1187),
            data_im_in => first_stage_im_out(1187),
            re_multiplicator => "1110100101010101", --- -0.354187011719 + j-0.935180664062
            im_multiplicator => "1100010000100110",
            data_re_out => mul_re_out(1187),
            data_im_out => mul_im_out(1187)
        );

 
    UMUL_1188 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1188),
            data_im_in => first_stage_im_out(1188),
            re_multiplicator => "1110011000010001", --- -0.405212402344 + j-0.914184570312
            im_multiplicator => "1100010101111110",
            data_re_out => mul_re_out(1188),
            data_im_out => mul_im_out(1188)
        );

 
    UMUL_1189 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1189),
            data_im_in => first_stage_im_out(1189),
            re_multiplicator => "1110001011100000", --- -0.455078125 + j-0.890441894531
            im_multiplicator => "1100011100000011",
            data_re_out => mul_re_out(1189),
            data_im_out => mul_im_out(1189)
        );

 
    UMUL_1190 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1190),
            data_im_in => first_stage_im_out(1190),
            re_multiplicator => "1101111111000110", --- -0.503540039062 + j-0.863952636719
            im_multiplicator => "1100100010110101",
            data_re_out => mul_re_out(1190),
            data_im_out => mul_im_out(1190)
        );

 
    UMUL_1191 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1191),
            data_im_in => first_stage_im_out(1191),
            re_multiplicator => "1101110011000101", --- -0.550476074219 + j-0.834838867188
            im_multiplicator => "1100101010010010",
            data_re_out => mul_re_out(1191),
            data_im_out => mul_im_out(1191)
        );

 
    UMUL_1192 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1192),
            data_im_in => first_stage_im_out(1192),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(1192),
            data_im_out => mul_im_out(1192)
        );

 
    UMUL_1193 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1193),
            data_im_in => first_stage_im_out(1193),
            re_multiplicator => "1101011100011001", --- -0.639099121094 + j-0.769104003906
            im_multiplicator => "1100111011000111",
            data_re_out => mul_re_out(1193),
            data_im_out => mul_im_out(1193)
        );

 
    UMUL_1194 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1194),
            data_im_in => first_stage_im_out(1194),
            re_multiplicator => "1101010001110001", --- -0.680603027344 + j-0.732666015625
            im_multiplicator => "1101000100011100",
            data_re_out => mul_re_out(1194),
            data_im_out => mul_im_out(1194)
        );

 
    UMUL_1195 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1195),
            data_im_in => first_stage_im_out(1195),
            re_multiplicator => "1101000111101011", --- -0.720031738281 + j-0.693969726562
            im_multiplicator => "1101001110010110",
            data_re_out => mul_re_out(1195),
            data_im_out => mul_im_out(1195)
        );

 
    UMUL_1196 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1196),
            data_im_in => first_stage_im_out(1196),
            re_multiplicator => "1100111110001010", --- -0.757202148438 + j-0.653198242188
            im_multiplicator => "1101011000110010",
            data_re_out => mul_re_out(1196),
            data_im_out => mul_im_out(1196)
        );

 
    UMUL_1197 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1197),
            data_im_in => first_stage_im_out(1197),
            re_multiplicator => "1100110101001110", --- -0.792114257812 + j-0.610412597656
            im_multiplicator => "1101100011101111",
            data_re_out => mul_re_out(1197),
            data_im_out => mul_im_out(1197)
        );

 
    UMUL_1198 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1198),
            data_im_in => first_stage_im_out(1198),
            re_multiplicator => "1100101100111010", --- -0.824584960938 + j-0.565734863281
            im_multiplicator => "1101101111001011",
            data_re_out => mul_re_out(1198),
            data_im_out => mul_im_out(1198)
        );

 
    UMUL_1199 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1199),
            data_im_in => first_stage_im_out(1199),
            re_multiplicator => "1100100101001111", --- -0.854553222656 + j-0.519348144531
            im_multiplicator => "1101111011000011",
            data_re_out => mul_re_out(1199),
            data_im_out => mul_im_out(1199)
        );

 
    UMUL_1200 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1200),
            data_im_in => first_stage_im_out(1200),
            re_multiplicator => "1100011110001111", --- -0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(1200),
            data_im_out => mul_im_out(1200)
        );

 
    UMUL_1201 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1201),
            data_im_in => first_stage_im_out(1201),
            re_multiplicator => "1100010111111010", --- -0.906616210938 + j-0.421997070312
            im_multiplicator => "1110010011111110",
            data_re_out => mul_re_out(1201),
            data_im_out => mul_im_out(1201)
        );

 
    UMUL_1202 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1202),
            data_im_in => first_stage_im_out(1202),
            re_multiplicator => "1100010010010011", --- -0.928527832031 + j-0.371337890625
            im_multiplicator => "1110100000111100",
            data_re_out => mul_re_out(1202),
            data_im_out => mul_im_out(1202)
        );

 
    UMUL_1203 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1203),
            data_im_in => first_stage_im_out(1203),
            re_multiplicator => "1100001101011011", --- -0.947570800781 + j-0.319519042969
            im_multiplicator => "1110101110001101",
            data_re_out => mul_re_out(1203),
            data_im_out => mul_im_out(1203)
        );

 
    UMUL_1204 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1204),
            data_im_in => first_stage_im_out(1204),
            re_multiplicator => "1100001001010001", --- -0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(1204),
            data_im_out => mul_im_out(1204)
        );

 
    UMUL_1205 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1205),
            data_im_in => first_stage_im_out(1205),
            re_multiplicator => "1100000101111000", --- -0.97705078125 + j-0.213134765625
            im_multiplicator => "1111001001011100",
            data_re_out => mul_re_out(1205),
            data_im_out => mul_im_out(1205)
        );

 
    UMUL_1206 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1206),
            data_im_in => first_stage_im_out(1206),
            re_multiplicator => "1100000011010000", --- -0.9873046875 + j-0.158874511719
            im_multiplicator => "1111010111010101",
            data_re_out => mul_re_out(1206),
            data_im_out => mul_im_out(1206)
        );

 
    UMUL_1207 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1207),
            data_im_in => first_stage_im_out(1207),
            re_multiplicator => "1100000001011001", --- -0.994567871094 + j-0.104125976562
            im_multiplicator => "1111100101010110",
            data_re_out => mul_re_out(1207),
            data_im_out => mul_im_out(1207)
        );

 
    UMUL_1208 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1208),
            data_im_in => first_stage_im_out(1208),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(1208),
            data_im_out => mul_im_out(1208)
        );

 
    UMUL_1209 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1209),
            data_im_in => first_stage_im_out(1209),
            re_multiplicator => "1100000000000000", --- -1.0 + j0.00616455078125
            im_multiplicator => "0000000001100101",
            data_re_out => mul_re_out(1209),
            data_im_out => mul_im_out(1209)
        );

 
    UMUL_1210 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1210),
            data_im_in => first_stage_im_out(1210),
            re_multiplicator => "1100000000011111", --- -0.998107910156 + j0.0613403320312
            im_multiplicator => "0000001111101101",
            data_re_out => mul_re_out(1210),
            data_im_out => mul_im_out(1210)
        );

 
    UMUL_1211 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1211),
            data_im_in => first_stage_im_out(1211),
            re_multiplicator => "1100000001101111", --- -0.993225097656 + j0.116333007812
            im_multiplicator => "0000011101110010",
            data_re_out => mul_re_out(1211),
            data_im_out => mul_im_out(1211)
        );

 
    UMUL_1212 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1212),
            data_im_in => first_stage_im_out(1212),
            re_multiplicator => "1100000011110001", --- -0.985290527344 + j0.170959472656
            im_multiplicator => "0000101011110001",
            data_re_out => mul_re_out(1212),
            data_im_out => mul_im_out(1212)
        );

 
    UMUL_1213 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1213),
            data_im_in => first_stage_im_out(1213),
            re_multiplicator => "1100000110100100", --- -0.974365234375 + j0.22509765625
            im_multiplicator => "0000111001101000",
            data_re_out => mul_re_out(1213),
            data_im_out => mul_im_out(1213)
        );

 
    UMUL_1214 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1214),
            data_im_in => first_stage_im_out(1214),
            re_multiplicator => "1100001010001000", --- -0.96044921875 + j0.278503417969
            im_multiplicator => "0001000111010011",
            data_re_out => mul_re_out(1214),
            data_im_out => mul_im_out(1214)
        );

 
    UMUL_1215 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1215),
            data_im_in => first_stage_im_out(1215),
            re_multiplicator => "1100001110011100", --- -0.943603515625 + j0.331115722656
            im_multiplicator => "0001010100110001",
            data_re_out => mul_re_out(1215),
            data_im_out => mul_im_out(1215)
        );

 
    UMUL_1216 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1216),
            data_im_in => first_stage_im_out(1216),
            data_re_out => mul_re_out(1216),
            data_im_out => mul_im_out(1216)
        );

 
    UMUL_1217 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1217),
            data_im_in => first_stage_im_out(1217),
            re_multiplicator => "0011111111100100", --- 0.998291015625 + j-0.0582885742188
            im_multiplicator => "1111110001000101",
            data_re_out => mul_re_out(1217),
            data_im_out => mul_im_out(1217)
        );

 
    UMUL_1218 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1218),
            data_im_in => first_stage_im_out(1218),
            re_multiplicator => "0011111110010001", --- 0.993225097656 + j-0.116333007812
            im_multiplicator => "1111100010001110",
            data_re_out => mul_re_out(1218),
            data_im_out => mul_im_out(1218)
        );

 
    UMUL_1219 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1219),
            data_im_in => first_stage_im_out(1219),
            re_multiplicator => "0011111100000110", --- 0.984741210938 + j-0.174011230469
            im_multiplicator => "1111010011011101",
            data_re_out => mul_re_out(1219),
            data_im_out => mul_im_out(1219)
        );

 
    UMUL_1220 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1220),
            data_im_in => first_stage_im_out(1220),
            re_multiplicator => "0011111001000101", --- 0.972961425781 + j-0.231079101562
            im_multiplicator => "1111000100110110",
            data_re_out => mul_re_out(1220),
            data_im_out => mul_im_out(1220)
        );

 
    UMUL_1221 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1221),
            data_im_in => first_stage_im_out(1221),
            re_multiplicator => "0011110101001101", --- 0.957824707031 + j-0.287353515625
            im_multiplicator => "1110110110011100",
            data_re_out => mul_re_out(1221),
            data_im_out => mul_im_out(1221)
        );

 
    UMUL_1222 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1222),
            data_im_in => first_stage_im_out(1222),
            re_multiplicator => "0011110000100000", --- 0.939453125 + j-0.342651367188
            im_multiplicator => "1110101000010010",
            data_re_out => mul_re_out(1222),
            data_im_out => mul_im_out(1222)
        );

 
    UMUL_1223 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1223),
            data_im_in => first_stage_im_out(1223),
            re_multiplicator => "0011101010111111", --- 0.917907714844 + j-0.396789550781
            im_multiplicator => "1110011010011011",
            data_re_out => mul_re_out(1223),
            data_im_out => mul_im_out(1223)
        );

 
    UMUL_1224 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1224),
            data_im_in => first_stage_im_out(1224),
            re_multiplicator => "0011100100101011", --- 0.893249511719 + j-0.449584960938
            im_multiplicator => "1110001100111010",
            data_re_out => mul_re_out(1224),
            data_im_out => mul_im_out(1224)
        );

 
    UMUL_1225 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1225),
            data_im_in => first_stage_im_out(1225),
            re_multiplicator => "0011011101100101", --- 0.865539550781 + j-0.500915527344
            im_multiplicator => "1101111111110001",
            data_re_out => mul_re_out(1225),
            data_im_out => mul_im_out(1225)
        );

 
    UMUL_1226 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1226),
            data_im_in => first_stage_im_out(1226),
            re_multiplicator => "0011010101101110", --- 0.834838867188 + j-0.550476074219
            im_multiplicator => "1101110011000101",
            data_re_out => mul_re_out(1226),
            data_im_out => mul_im_out(1226)
        );

 
    UMUL_1227 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1227),
            data_im_in => first_stage_im_out(1227),
            re_multiplicator => "0011001101001010", --- 0.801391601562 + j-0.59814453125
            im_multiplicator => "1101100110111000",
            data_re_out => mul_re_out(1227),
            data_im_out => mul_im_out(1227)
        );

 
    UMUL_1228 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1228),
            data_im_in => first_stage_im_out(1228),
            re_multiplicator => "0011000011111001", --- 0.765197753906 + j-0.643859863281
            im_multiplicator => "1101011011001011",
            data_re_out => mul_re_out(1228),
            data_im_out => mul_im_out(1228)
        );

 
    UMUL_1229 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1229),
            data_im_in => first_stage_im_out(1229),
            re_multiplicator => "0010111001111101", --- 0.726379394531 + j-0.687316894531
            im_multiplicator => "1101010000000011",
            data_re_out => mul_re_out(1229),
            data_im_out => mul_im_out(1229)
        );

 
    UMUL_1230 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1230),
            data_im_in => first_stage_im_out(1230),
            re_multiplicator => "0010101111011000", --- 0.68505859375 + j-0.728454589844
            im_multiplicator => "1101000101100001",
            data_re_out => mul_re_out(1230),
            data_im_out => mul_im_out(1230)
        );

 
    UMUL_1231 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1231),
            data_im_in => first_stage_im_out(1231),
            re_multiplicator => "0010100100001110", --- 0.641479492188 + j-0.767150878906
            im_multiplicator => "1100111011100111",
            data_re_out => mul_re_out(1231),
            data_im_out => mul_im_out(1231)
        );

 
    UMUL_1232 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1232),
            data_im_in => first_stage_im_out(1232),
            re_multiplicator => "0010011000100000", --- 0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(1232),
            data_im_out => mul_im_out(1232)
        );

 
    UMUL_1233 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1233),
            data_im_in => first_stage_im_out(1233),
            re_multiplicator => "0010001100010001", --- 0.547912597656 + j-0.836547851562
            im_multiplicator => "1100101001110110",
            data_re_out => mul_re_out(1233),
            data_im_out => mul_im_out(1233)
        );

 
    UMUL_1234 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1234),
            data_im_in => first_stage_im_out(1234),
            re_multiplicator => "0001111111100011", --- 0.498229980469 + j-0.867065429688
            im_multiplicator => "1100100010000010",
            data_re_out => mul_re_out(1234),
            data_im_out => mul_im_out(1234)
        );

 
    UMUL_1235 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1235),
            data_im_in => first_stage_im_out(1235),
            re_multiplicator => "0001110010011001", --- 0.446838378906 + j-0.894592285156
            im_multiplicator => "1100011010111111",
            data_re_out => mul_re_out(1235),
            data_im_out => mul_im_out(1235)
        );

 
    UMUL_1236 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1236),
            data_im_in => first_stage_im_out(1236),
            re_multiplicator => "0001100100110111", --- 0.393981933594 + j-0.919128417969
            im_multiplicator => "1100010100101101",
            data_re_out => mul_re_out(1236),
            data_im_out => mul_im_out(1236)
        );

 
    UMUL_1237 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1237),
            data_im_in => first_stage_im_out(1237),
            re_multiplicator => "0001010110111111", --- 0.339782714844 + j-0.940490722656
            im_multiplicator => "1100001111001111",
            data_re_out => mul_re_out(1237),
            data_im_out => mul_im_out(1237)
        );

 
    UMUL_1238 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1238),
            data_im_in => first_stage_im_out(1238),
            re_multiplicator => "0001001000110100", --- 0.284423828125 + j-0.958679199219
            im_multiplicator => "1100001010100101",
            data_re_out => mul_re_out(1238),
            data_im_out => mul_im_out(1238)
        );

 
    UMUL_1239 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1239),
            data_im_in => first_stage_im_out(1239),
            re_multiplicator => "0000111010011001", --- 0.228088378906 + j-0.9736328125
            im_multiplicator => "1100000110110000",
            data_re_out => mul_re_out(1239),
            data_im_out => mul_im_out(1239)
        );

 
    UMUL_1240 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1240),
            data_im_in => first_stage_im_out(1240),
            re_multiplicator => "0000101011110001", --- 0.170959472656 + j-0.985290527344
            im_multiplicator => "1100000011110001",
            data_re_out => mul_re_out(1240),
            data_im_out => mul_im_out(1240)
        );

 
    UMUL_1241 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1241),
            data_im_in => first_stage_im_out(1241),
            re_multiplicator => "0000011101000000", --- 0.11328125 + j-0.993591308594
            im_multiplicator => "1100000001101001",
            data_re_out => mul_re_out(1241),
            data_im_out => mul_im_out(1241)
        );

 
    UMUL_1242 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1242),
            data_im_in => first_stage_im_out(1242),
            re_multiplicator => "0000001110001000", --- 0.05517578125 + j-0.998474121094
            im_multiplicator => "1100000000011001",
            data_re_out => mul_re_out(1242),
            data_im_out => mul_im_out(1242)
        );

 
    UMUL_1243 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1243),
            data_im_in => first_stage_im_out(1243),
            re_multiplicator => "1111111111001110", --- -0.0030517578125 + j-1.0
            im_multiplicator => "1100000000000000",
            data_re_out => mul_re_out(1243),
            data_im_out => mul_im_out(1243)
        );

 
    UMUL_1244 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1244),
            data_im_in => first_stage_im_out(1244),
            re_multiplicator => "1111110000010011", --- -0.0613403320312 + j-0.998107910156
            im_multiplicator => "1100000000011111",
            data_re_out => mul_re_out(1244),
            data_im_out => mul_im_out(1244)
        );

 
    UMUL_1245 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1245),
            data_im_in => first_stage_im_out(1245),
            re_multiplicator => "1111100001011100", --- -0.119384765625 + j-0.992858886719
            im_multiplicator => "1100000001110101",
            data_re_out => mul_re_out(1245),
            data_im_out => mul_im_out(1245)
        );

 
    UMUL_1246 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1246),
            data_im_in => first_stage_im_out(1246),
            re_multiplicator => "1111010010101100", --- -0.177001953125 + j-0.984191894531
            im_multiplicator => "1100000100000011",
            data_re_out => mul_re_out(1246),
            data_im_out => mul_im_out(1246)
        );

 
    UMUL_1247 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1247),
            data_im_in => first_stage_im_out(1247),
            re_multiplicator => "1111000100000101", --- -0.234069824219 + j-0.972229003906
            im_multiplicator => "1100000111000111",
            data_re_out => mul_re_out(1247),
            data_im_out => mul_im_out(1247)
        );

 
    UMUL_1248 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1248),
            data_im_in => first_stage_im_out(1248),
            re_multiplicator => "1110110101101100", --- -0.290283203125 + j-0.956970214844
            im_multiplicator => "1100001011000001",
            data_re_out => mul_re_out(1248),
            data_im_out => mul_im_out(1248)
        );

 
    UMUL_1249 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1249),
            data_im_in => first_stage_im_out(1249),
            re_multiplicator => "1110100111100011", --- -0.345520019531 + j-0.938415527344
            im_multiplicator => "1100001111110001",
            data_re_out => mul_re_out(1249),
            data_im_out => mul_im_out(1249)
        );

 
    UMUL_1250 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1250),
            data_im_in => first_stage_im_out(1250),
            re_multiplicator => "1110011001101101", --- -0.399597167969 + j-0.916687011719
            im_multiplicator => "1100010101010101",
            data_re_out => mul_re_out(1250),
            data_im_out => mul_im_out(1250)
        );

 
    UMUL_1251 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1251),
            data_im_in => first_stage_im_out(1251),
            re_multiplicator => "1110001100001101", --- -0.452331542969 + j-0.891845703125
            im_multiplicator => "1100011011101100",
            data_re_out => mul_re_out(1251),
            data_im_out => mul_im_out(1251)
        );

 
    UMUL_1252 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1252),
            data_im_in => first_stage_im_out(1252),
            re_multiplicator => "1101111111000110", --- -0.503540039062 + j-0.863952636719
            im_multiplicator => "1100100010110101",
            data_re_out => mul_re_out(1252),
            data_im_out => mul_im_out(1252)
        );

 
    UMUL_1253 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1253),
            data_im_in => first_stage_im_out(1253),
            re_multiplicator => "1101110010011011", --- -0.553039550781 + j-0.833190917969
            im_multiplicator => "1100101010101101",
            data_re_out => mul_re_out(1253),
            data_im_out => mul_im_out(1253)
        );

 
    UMUL_1254 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1254),
            data_im_in => first_stage_im_out(1254),
            re_multiplicator => "1101100110001111", --- -0.600646972656 + j-0.799560546875
            im_multiplicator => "1100110011010100",
            data_re_out => mul_re_out(1254),
            data_im_out => mul_im_out(1254)
        );

 
    UMUL_1255 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1255),
            data_im_in => first_stage_im_out(1255),
            re_multiplicator => "1101011010100101", --- -0.646179199219 + j-0.76318359375
            im_multiplicator => "1100111100101000",
            data_re_out => mul_re_out(1255),
            data_im_out => mul_im_out(1255)
        );

 
    UMUL_1256 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1256),
            data_im_in => first_stage_im_out(1256),
            re_multiplicator => "1101001111011111", --- -0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(1256),
            data_im_out => mul_im_out(1256)
        );

 
    UMUL_1257 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1257),
            data_im_in => first_stage_im_out(1257),
            re_multiplicator => "1101000100111110", --- -0.730590820312 + j-0.682861328125
            im_multiplicator => "1101010001001100",
            data_re_out => mul_re_out(1257),
            data_im_out => mul_im_out(1257)
        );

 
    UMUL_1258 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1258),
            data_im_in => first_stage_im_out(1258),
            re_multiplicator => "1100111011000111", --- -0.769104003906 + j-0.639099121094
            im_multiplicator => "1101011100011001",
            data_re_out => mul_re_out(1258),
            data_im_out => mul_im_out(1258)
        );

 
    UMUL_1259 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1259),
            data_im_in => first_stage_im_out(1259),
            re_multiplicator => "1100110001111010", --- -0.805053710938 + j-0.59326171875
            im_multiplicator => "1101101000001000",
            data_re_out => mul_re_out(1259),
            data_im_out => mul_im_out(1259)
        );

 
    UMUL_1260 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1260),
            data_im_in => first_stage_im_out(1260),
            re_multiplicator => "1100101001011011", --- -0.838195800781 + j-0.545349121094
            im_multiplicator => "1101110100011001",
            data_re_out => mul_re_out(1260),
            data_im_out => mul_im_out(1260)
        );

 
    UMUL_1261 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1261),
            data_im_in => first_stage_im_out(1261),
            re_multiplicator => "1100100001101001", --- -0.868591308594 + j-0.495544433594
            im_multiplicator => "1110000001001001",
            data_re_out => mul_re_out(1261),
            data_im_out => mul_im_out(1261)
        );

 
    UMUL_1262 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1262),
            data_im_in => first_stage_im_out(1262),
            re_multiplicator => "1100011010101000", --- -0.89599609375 + j-0.444091796875
            im_multiplicator => "1110001110010100",
            data_re_out => mul_re_out(1262),
            data_im_out => mul_im_out(1262)
        );

 
    UMUL_1263 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1263),
            data_im_in => first_stage_im_out(1263),
            re_multiplicator => "1100010100011010", --- -0.920288085938 + j-0.391174316406
            im_multiplicator => "1110011011110111",
            data_re_out => mul_re_out(1263),
            data_im_out => mul_im_out(1263)
        );

 
    UMUL_1264 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1264),
            data_im_in => first_stage_im_out(1264),
            re_multiplicator => "1100001110111110", --- -0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(1264),
            data_im_out => mul_im_out(1264)
        );

 
    UMUL_1265 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1265),
            data_im_in => first_stage_im_out(1265),
            re_multiplicator => "1100001010010110", --- -0.959594726562 + j-0.281494140625
            im_multiplicator => "1110110111111100",
            data_re_out => mul_re_out(1265),
            data_im_out => mul_im_out(1265)
        );

 
    UMUL_1266 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1266),
            data_im_in => first_stage_im_out(1266),
            re_multiplicator => "1100000110100100", --- -0.974365234375 + j-0.22509765625
            im_multiplicator => "1111000110011000",
            data_re_out => mul_re_out(1266),
            data_im_out => mul_im_out(1266)
        );

 
    UMUL_1267 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1267),
            data_im_in => first_stage_im_out(1267),
            re_multiplicator => "1100000011101001", --- -0.985778808594 + j-0.16796875
            im_multiplicator => "1111010101000000",
            data_re_out => mul_re_out(1267),
            data_im_out => mul_im_out(1267)
        );

 
    UMUL_1268 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1268),
            data_im_in => first_stage_im_out(1268),
            re_multiplicator => "1100000001100100", --- -0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(1268),
            data_im_out => mul_im_out(1268)
        );

 
    UMUL_1269 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1269),
            data_im_in => first_stage_im_out(1269),
            re_multiplicator => "1100000000010110", --- -0.998657226562 + j-0.0521240234375
            im_multiplicator => "1111110010101010",
            data_re_out => mul_re_out(1269),
            data_im_out => mul_im_out(1269)
        );

 
    UMUL_1270 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1270),
            data_im_in => first_stage_im_out(1270),
            re_multiplicator => "1100000000000000", --- -1.0 + j0.00616455078125
            im_multiplicator => "0000000001100101",
            data_re_out => mul_re_out(1270),
            data_im_out => mul_im_out(1270)
        );

 
    UMUL_1271 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1271),
            data_im_in => first_stage_im_out(1271),
            re_multiplicator => "1100000000100010", --- -0.997924804688 + j0.0643920898438
            im_multiplicator => "0000010000011111",
            data_re_out => mul_re_out(1271),
            data_im_out => mul_im_out(1271)
        );

 
    UMUL_1272 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1272),
            data_im_in => first_stage_im_out(1272),
            re_multiplicator => "1100000001111011", --- -0.992492675781 + j0.122436523438
            im_multiplicator => "0000011111010110",
            data_re_out => mul_re_out(1272),
            data_im_out => mul_im_out(1272)
        );

 
    UMUL_1273 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1273),
            data_im_in => first_stage_im_out(1273),
            re_multiplicator => "1100000100001100", --- -0.983642578125 + j0.179992675781
            im_multiplicator => "0000101110000101",
            data_re_out => mul_re_out(1273),
            data_im_out => mul_im_out(1273)
        );

 
    UMUL_1274 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1274),
            data_im_in => first_stage_im_out(1274),
            re_multiplicator => "1100000111010011", --- -0.971496582031 + j0.236999511719
            im_multiplicator => "0000111100101011",
            data_re_out => mul_re_out(1274),
            data_im_out => mul_im_out(1274)
        );

 
    UMUL_1275 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1275),
            data_im_in => first_stage_im_out(1275),
            re_multiplicator => "1100001011010000", --- -0.9560546875 + j0.293212890625
            im_multiplicator => "0001001011000100",
            data_re_out => mul_re_out(1275),
            data_im_out => mul_im_out(1275)
        );

 
    UMUL_1276 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1276),
            data_im_in => first_stage_im_out(1276),
            re_multiplicator => "1100010000000011", --- -0.937316894531 + j0.348388671875
            im_multiplicator => "0001011001001100",
            data_re_out => mul_re_out(1276),
            data_im_out => mul_im_out(1276)
        );

 
    UMUL_1277 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1277),
            data_im_in => first_stage_im_out(1277),
            re_multiplicator => "1100010101101001", --- -0.915466308594 + j0.402404785156
            im_multiplicator => "0001100111000001",
            data_re_out => mul_re_out(1277),
            data_im_out => mul_im_out(1277)
        );

 
    UMUL_1278 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1278),
            data_im_in => first_stage_im_out(1278),
            re_multiplicator => "1100011100000011", --- -0.890441894531 + j0.455078125
            im_multiplicator => "0001110100100000",
            data_re_out => mul_re_out(1278),
            data_im_out => mul_im_out(1278)
        );

 
    UMUL_1279 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1279),
            data_im_in => first_stage_im_out(1279),
            re_multiplicator => "1100100011001110", --- -0.862426757812 + j0.506164550781
            im_multiplicator => "0010000001100101",
            data_re_out => mul_re_out(1279),
            data_im_out => mul_im_out(1279)
        );

 
    UMUL_1280 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1280),
            data_im_in => first_stage_im_out(1280),
            data_re_out => mul_re_out(1280),
            data_im_out => mul_im_out(1280)
        );

 
    UMUL_1281 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1281),
            data_im_in => first_stage_im_out(1281),
            re_multiplicator => "0011111111100001", --- 0.998107910156 + j-0.0613403320312
            im_multiplicator => "1111110000010011",
            data_re_out => mul_re_out(1281),
            data_im_out => mul_im_out(1281)
        );

 
    UMUL_1282 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1282),
            data_im_in => first_stage_im_out(1282),
            re_multiplicator => "0011111110000101", --- 0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(1282),
            data_im_out => mul_im_out(1282)
        );

 
    UMUL_1283 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1283),
            data_im_in => first_stage_im_out(1283),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(1283),
            data_im_out => mul_im_out(1283)
        );

 
    UMUL_1284 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1284),
            data_im_in => first_stage_im_out(1284),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(1284),
            data_im_out => mul_im_out(1284)
        );

 
    UMUL_1285 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1285),
            data_im_in => first_stage_im_out(1285),
            re_multiplicator => "0011110100000011", --- 0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(1285),
            data_im_out => mul_im_out(1285)
        );

 
    UMUL_1286 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1286),
            data_im_in => first_stage_im_out(1286),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(1286),
            data_im_out => mul_im_out(1286)
        );

 
    UMUL_1287 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1287),
            data_im_in => first_stage_im_out(1287),
            re_multiplicator => "0011101000110000", --- 0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(1287),
            data_im_out => mul_im_out(1287)
        );

 
    UMUL_1288 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1288),
            data_im_in => first_stage_im_out(1288),
            re_multiplicator => "0011100001110001", --- 0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(1288),
            data_im_out => mul_im_out(1288)
        );

 
    UMUL_1289 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1289),
            data_im_in => first_stage_im_out(1289),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(1289),
            data_im_out => mul_im_out(1289)
        );

 
    UMUL_1290 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1290),
            data_im_in => first_stage_im_out(1290),
            re_multiplicator => "0011010001010011", --- 0.817565917969 + j-0.575805664062
            im_multiplicator => "1101101100100110",
            data_re_out => mul_re_out(1290),
            data_im_out => mul_im_out(1290)
        );

 
    UMUL_1291 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1291),
            data_im_in => first_stage_im_out(1291),
            re_multiplicator => "0011000111111000", --- 0.78076171875 + j-0.624877929688
            im_multiplicator => "1101100000000010",
            data_re_out => mul_re_out(1291),
            data_im_out => mul_im_out(1291)
        );

 
    UMUL_1292 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1292),
            data_im_in => first_stage_im_out(1292),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(1292),
            data_im_out => mul_im_out(1292)
        );

 
    UMUL_1293 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1293),
            data_im_in => first_stage_im_out(1293),
            re_multiplicator => "0010110010110010", --- 0.698364257812 + j-0.715759277344
            im_multiplicator => "1101001000110001",
            data_re_out => mul_re_out(1293),
            data_im_out => mul_im_out(1293)
        );

 
    UMUL_1294 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1294),
            data_im_in => first_stage_im_out(1294),
            re_multiplicator => "0010100111001110", --- 0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(1294),
            data_im_out => mul_im_out(1294)
        );

 
    UMUL_1295 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1295),
            data_im_in => first_stage_im_out(1295),
            re_multiplicator => "0010011011000001", --- 0.605529785156 + j-0.795837402344
            im_multiplicator => "1100110100010001",
            data_re_out => mul_re_out(1295),
            data_im_out => mul_im_out(1295)
        );

 
    UMUL_1296 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1296),
            data_im_in => first_stage_im_out(1296),
            re_multiplicator => "0010001110001110", --- 0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(1296),
            data_im_out => mul_im_out(1296)
        );

 
    UMUL_1297 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1297),
            data_im_in => first_stage_im_out(1297),
            re_multiplicator => "0010000000111010", --- 0.503540039062 + j-0.863952636719
            im_multiplicator => "1100100010110101",
            data_re_out => mul_re_out(1297),
            data_im_out => mul_im_out(1297)
        );

 
    UMUL_1298 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1298),
            data_im_in => first_stage_im_out(1298),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(1298),
            data_im_out => mul_im_out(1298)
        );

 
    UMUL_1299 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1299),
            data_im_in => first_stage_im_out(1299),
            re_multiplicator => "0001100100110111", --- 0.393981933594 + j-0.919128417969
            im_multiplicator => "1100010100101101",
            data_re_out => mul_re_out(1299),
            data_im_out => mul_im_out(1299)
        );

 
    UMUL_1300 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1300),
            data_im_in => first_stage_im_out(1300),
            re_multiplicator => "0001010110010000", --- 0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(1300),
            data_im_out => mul_im_out(1300)
        );

 
    UMUL_1301 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1301),
            data_im_in => first_stage_im_out(1301),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(1301),
            data_im_out => mul_im_out(1301)
        );

 
    UMUL_1302 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1302),
            data_im_in => first_stage_im_out(1302),
            re_multiplicator => "0000111000000110", --- 0.219116210938 + j-0.975708007812
            im_multiplicator => "1100000110001110",
            data_re_out => mul_re_out(1302),
            data_im_out => mul_im_out(1302)
        );

 
    UMUL_1303 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1303),
            data_im_in => first_stage_im_out(1303),
            re_multiplicator => "0000101000101011", --- 0.158874511719 + j-0.9873046875
            im_multiplicator => "1100000011010000",
            data_re_out => mul_re_out(1303),
            data_im_out => mul_im_out(1303)
        );

 
    UMUL_1304 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1304),
            data_im_in => first_stage_im_out(1304),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(1304),
            data_im_out => mul_im_out(1304)
        );

 
    UMUL_1305 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1305),
            data_im_in => first_stage_im_out(1305),
            re_multiplicator => "0000001001011011", --- 0.0368041992188 + j-0.999328613281
            im_multiplicator => "1100000000001011",
            data_re_out => mul_re_out(1305),
            data_im_out => mul_im_out(1305)
        );

 
    UMUL_1306 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1306),
            data_im_in => first_stage_im_out(1306),
            re_multiplicator => "1111111001101110", --- -0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(1306),
            data_im_out => mul_im_out(1306)
        );

 
    UMUL_1307 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1307),
            data_im_in => first_stage_im_out(1307),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(1307),
            data_im_out => mul_im_out(1307)
        );

 
    UMUL_1308 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1308),
            data_im_in => first_stage_im_out(1308),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(1308),
            data_im_out => mul_im_out(1308)
        );

 
    UMUL_1309 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1309),
            data_im_in => first_stage_im_out(1309),
            re_multiplicator => "1111001010111111", --- -0.207092285156 + j-0.978332519531
            im_multiplicator => "1100000101100011",
            data_re_out => mul_re_out(1309),
            data_im_out => mul_im_out(1309)
        );

 
    UMUL_1310 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1310),
            data_im_in => first_stage_im_out(1310),
            re_multiplicator => "1110111011101110", --- -0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(1310),
            data_im_out => mul_im_out(1310)
        );

 
    UMUL_1311 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1311),
            data_im_in => first_stage_im_out(1311),
            re_multiplicator => "1110101100101110", --- -0.325317382812 + j-0.945617675781
            im_multiplicator => "1100001101111011",
            data_re_out => mul_re_out(1311),
            data_im_out => mul_im_out(1311)
        );

 
    UMUL_1312 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1312),
            data_im_in => first_stage_im_out(1312),
            re_multiplicator => "1110011110000010", --- -0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(1312),
            data_im_out => mul_im_out(1312)
        );

 
    UMUL_1313 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1313),
            data_im_in => first_stage_im_out(1313),
            re_multiplicator => "1110001111101110", --- -0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(1313),
            data_im_out => mul_im_out(1313)
        );

 
    UMUL_1314 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1314),
            data_im_in => first_stage_im_out(1314),
            re_multiplicator => "1110000001110100", --- -0.492919921875 + j-0.8701171875
            im_multiplicator => "1100100001010000",
            data_re_out => mul_re_out(1314),
            data_im_out => mul_im_out(1314)
        );

 
    UMUL_1315 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1315),
            data_im_in => first_stage_im_out(1315),
            re_multiplicator => "1101110100011001", --- -0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(1315),
            data_im_out => mul_im_out(1315)
        );

 
    UMUL_1316 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1316),
            data_im_in => first_stage_im_out(1316),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(1316),
            data_im_out => mul_im_out(1316)
        );

 
    UMUL_1317 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1317),
            data_im_in => first_stage_im_out(1317),
            re_multiplicator => "1101011011001011", --- -0.643859863281 + j-0.765197753906
            im_multiplicator => "1100111100000111",
            data_re_out => mul_re_out(1317),
            data_im_out => mul_im_out(1317)
        );

 
    UMUL_1318 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1318),
            data_im_in => first_stage_im_out(1318),
            re_multiplicator => "1101001111011111", --- -0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(1318),
            data_im_out => mul_im_out(1318)
        );

 
    UMUL_1319 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1319),
            data_im_in => first_stage_im_out(1319),
            re_multiplicator => "1101000100011100", --- -0.732666015625 + j-0.680603027344
            im_multiplicator => "1101010001110001",
            data_re_out => mul_re_out(1319),
            data_im_out => mul_im_out(1319)
        );

 
    UMUL_1320 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1320),
            data_im_in => first_stage_im_out(1320),
            re_multiplicator => "1100111010000111", --- -0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(1320),
            data_im_out => mul_im_out(1320)
        );

 
    UMUL_1321 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1321),
            data_im_in => first_stage_im_out(1321),
            re_multiplicator => "1100110000100001", --- -0.810485839844 + j-0.585815429688
            im_multiplicator => "1101101010000010",
            data_re_out => mul_re_out(1321),
            data_im_out => mul_im_out(1321)
        );

 
    UMUL_1322 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1322),
            data_im_in => first_stage_im_out(1322),
            re_multiplicator => "1100100111101110", --- -0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(1322),
            data_im_out => mul_im_out(1322)
        );

 
    UMUL_1323 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1323),
            data_im_in => first_stage_im_out(1323),
            re_multiplicator => "1100011111101110", --- -0.876098632812 + j-0.482177734375
            im_multiplicator => "1110000100100100",
            data_re_out => mul_re_out(1323),
            data_im_out => mul_im_out(1323)
        );

 
    UMUL_1324 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1324),
            data_im_in => first_stage_im_out(1324),
            re_multiplicator => "1100011000100101", --- -0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(1324),
            data_im_out => mul_im_out(1324)
        );

 
    UMUL_1325 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1325),
            data_im_in => first_stage_im_out(1325),
            re_multiplicator => "1100010010010011", --- -0.928527832031 + j-0.371337890625
            im_multiplicator => "1110100000111100",
            data_re_out => mul_re_out(1325),
            data_im_out => mul_im_out(1325)
        );

 
    UMUL_1326 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1326),
            data_im_in => first_stage_im_out(1326),
            re_multiplicator => "1100001100111011", --- -0.949523925781 + j-0.313659667969
            im_multiplicator => "1110101111101101",
            data_re_out => mul_re_out(1326),
            data_im_out => mul_im_out(1326)
        );

 
    UMUL_1327 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1327),
            data_im_in => first_stage_im_out(1327),
            re_multiplicator => "1100001000011101", --- -0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(1327),
            data_im_out => mul_im_out(1327)
        );

 
    UMUL_1328 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1328),
            data_im_in => first_stage_im_out(1328),
            re_multiplicator => "1100000100111011", --- -0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(1328),
            data_im_out => mul_im_out(1328)
        );

 
    UMUL_1329 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1329),
            data_im_in => first_stage_im_out(1329),
            re_multiplicator => "1100000010010101", --- -0.990905761719 + j-0.134582519531
            im_multiplicator => "1111011101100011",
            data_re_out => mul_re_out(1329),
            data_im_out => mul_im_out(1329)
        );

 
    UMUL_1330 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1330),
            data_im_in => first_stage_im_out(1330),
            re_multiplicator => "1100000000101100", --- -0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(1330),
            data_im_out => mul_im_out(1330)
        );

 
    UMUL_1331 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1331),
            data_im_in => first_stage_im_out(1331),
            re_multiplicator => "1100000000000001", --- -0.999938964844 + j-0.0122680664062
            im_multiplicator => "1111111100110111",
            data_re_out => mul_re_out(1331),
            data_im_out => mul_im_out(1331)
        );

 
    UMUL_1332 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1332),
            data_im_in => first_stage_im_out(1332),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j0.049072265625
            im_multiplicator => "0000001100100100",
            data_re_out => mul_re_out(1332),
            data_im_out => mul_im_out(1332)
        );

 
    UMUL_1333 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1333),
            data_im_in => first_stage_im_out(1333),
            re_multiplicator => "1100000001100100", --- -0.993896484375 + j0.110229492188
            im_multiplicator => "0000011100001110",
            data_re_out => mul_re_out(1333),
            data_im_out => mul_im_out(1333)
        );

 
    UMUL_1334 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1334),
            data_im_in => first_stage_im_out(1334),
            re_multiplicator => "1100000011110001", --- -0.985290527344 + j0.170959472656
            im_multiplicator => "0000101011110001",
            data_re_out => mul_re_out(1334),
            data_im_out => mul_im_out(1334)
        );

 
    UMUL_1335 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1335),
            data_im_in => first_stage_im_out(1335),
            re_multiplicator => "1100000110111011", --- -0.972961425781 + j0.231079101562
            im_multiplicator => "0000111011001010",
            data_re_out => mul_re_out(1335),
            data_im_out => mul_im_out(1335)
        );

 
    UMUL_1336 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1336),
            data_im_in => first_stage_im_out(1336),
            re_multiplicator => "1100001011000001", --- -0.956970214844 + j0.290283203125
            im_multiplicator => "0001001010010100",
            data_re_out => mul_re_out(1336),
            data_im_out => mul_im_out(1336)
        );

 
    UMUL_1337 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1337),
            data_im_in => first_stage_im_out(1337),
            re_multiplicator => "1100010000000011", --- -0.937316894531 + j0.348388671875
            im_multiplicator => "0001011001001100",
            data_re_out => mul_re_out(1337),
            data_im_out => mul_im_out(1337)
        );

 
    UMUL_1338 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1338),
            data_im_in => first_stage_im_out(1338),
            re_multiplicator => "1100010101111110", --- -0.914184570312 + j0.405212402344
            im_multiplicator => "0001100111101111",
            data_re_out => mul_re_out(1338),
            data_im_out => mul_im_out(1338)
        );

 
    UMUL_1339 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1339),
            data_im_in => first_stage_im_out(1339),
            re_multiplicator => "1100011100110001", --- -0.887634277344 + j0.460510253906
            im_multiplicator => "0001110101111001",
            data_re_out => mul_re_out(1339),
            data_im_out => mul_im_out(1339)
        );

 
    UMUL_1340 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1340),
            data_im_in => first_stage_im_out(1340),
            re_multiplicator => "1100100100011011", --- -0.857727050781 + j0.514099121094
            im_multiplicator => "0010000011100111",
            data_re_out => mul_re_out(1340),
            data_im_out => mul_im_out(1340)
        );

 
    UMUL_1341 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1341),
            data_im_in => first_stage_im_out(1341),
            re_multiplicator => "1100101100111010", --- -0.824584960938 + j0.565734863281
            im_multiplicator => "0010010000110101",
            data_re_out => mul_re_out(1341),
            data_im_out => mul_im_out(1341)
        );

 
    UMUL_1342 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1342),
            data_im_in => first_stage_im_out(1342),
            re_multiplicator => "1100110110001100", --- -0.788330078125 + j0.615234375
            im_multiplicator => "0010011101100000",
            data_re_out => mul_re_out(1342),
            data_im_out => mul_im_out(1342)
        );

 
    UMUL_1343 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1343),
            data_im_in => first_stage_im_out(1343),
            re_multiplicator => "1101000000001110", --- -0.749145507812 + j0.662414550781
            im_multiplicator => "0010101001100101",
            data_re_out => mul_re_out(1343),
            data_im_out => mul_im_out(1343)
        );

 
    UMUL_1344 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1344),
            data_im_in => first_stage_im_out(1344),
            data_re_out => mul_re_out(1344),
            data_im_out => mul_im_out(1344)
        );

 
    UMUL_1345 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1345),
            data_im_in => first_stage_im_out(1345),
            re_multiplicator => "0011111111011110", --- 0.997924804688 + j-0.0643920898438
            im_multiplicator => "1111101111100001",
            data_re_out => mul_re_out(1345),
            data_im_out => mul_im_out(1345)
        );

 
    UMUL_1346 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1346),
            data_im_in => first_stage_im_out(1346),
            re_multiplicator => "0011111101111000", --- 0.99169921875 + j-0.128479003906
            im_multiplicator => "1111011111000111",
            data_re_out => mul_re_out(1346),
            data_im_out => mul_im_out(1346)
        );

 
    UMUL_1347 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1347),
            data_im_in => first_stage_im_out(1347),
            re_multiplicator => "0011111011001111", --- 0.981384277344 + j-0.192077636719
            im_multiplicator => "1111001110110101",
            data_re_out => mul_re_out(1347),
            data_im_out => mul_im_out(1347)
        );

 
    UMUL_1348 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1348),
            data_im_in => first_stage_im_out(1348),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(1348),
            data_im_out => mul_im_out(1348)
        );

 
    UMUL_1349 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1349),
            data_im_in => first_stage_im_out(1349),
            re_multiplicator => "0011110010110101", --- 0.948547363281 + j-0.316589355469
            im_multiplicator => "1110101110111101",
            data_re_out => mul_re_out(1349),
            data_im_out => mul_im_out(1349)
        );

 
    UMUL_1350 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1350),
            data_im_in => first_stage_im_out(1350),
            re_multiplicator => "0011101101000111", --- 0.926208496094 + j-0.377014160156
            im_multiplicator => "1110011111011111",
            data_re_out => mul_re_out(1350),
            data_im_out => mul_im_out(1350)
        );

 
    UMUL_1351 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1351),
            data_im_in => first_stage_im_out(1351),
            re_multiplicator => "0011100110011010", --- 0.900024414062 + j-0.435852050781
            im_multiplicator => "1110010000011011",
            data_re_out => mul_re_out(1351),
            data_im_out => mul_im_out(1351)
        );

 
    UMUL_1352 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1352),
            data_im_in => first_stage_im_out(1352),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(1352),
            data_im_out => mul_im_out(1352)
        );

 
    UMUL_1353 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1353),
            data_im_in => first_stage_im_out(1353),
            re_multiplicator => "0011010110001010", --- 0.836547851562 + j-0.547912597656
            im_multiplicator => "1101110011101111",
            data_re_out => mul_re_out(1353),
            data_im_out => mul_im_out(1353)
        );

 
    UMUL_1354 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1354),
            data_im_in => first_stage_im_out(1354),
            re_multiplicator => "0011001100101100", --- 0.799560546875 + j-0.600646972656
            im_multiplicator => "1101100110001111",
            data_re_out => mul_re_out(1354),
            data_im_out => mul_im_out(1354)
        );

 
    UMUL_1355 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1355),
            data_im_in => first_stage_im_out(1355),
            re_multiplicator => "0011000010010111", --- 0.759216308594 + j-0.650817871094
            im_multiplicator => "1101011001011001",
            data_re_out => mul_re_out(1355),
            data_im_out => mul_im_out(1355)
        );

 
    UMUL_1356 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1356),
            data_im_in => first_stage_im_out(1356),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(1356),
            data_im_out => mul_im_out(1356)
        );

 
    UMUL_1357 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1357),
            data_im_in => first_stage_im_out(1357),
            re_multiplicator => "0010101011010110", --- 0.669311523438 + j-0.742980957031
            im_multiplicator => "1101000001110011",
            data_re_out => mul_re_out(1357),
            data_im_out => mul_im_out(1357)
        );

 
    UMUL_1358 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1358),
            data_im_in => first_stage_im_out(1358),
            re_multiplicator => "0010011110101111", --- 0.620056152344 + j-0.784545898438
            im_multiplicator => "1100110111001010",
            data_re_out => mul_re_out(1358),
            data_im_out => mul_im_out(1358)
        );

 
    UMUL_1359 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1359),
            data_im_in => first_stage_im_out(1359),
            re_multiplicator => "0010010001011110", --- 0.568237304688 + j-0.822875976562
            im_multiplicator => "1100101101010110",
            data_re_out => mul_re_out(1359),
            data_im_out => mul_im_out(1359)
        );

 
    UMUL_1360 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1360),
            data_im_in => first_stage_im_out(1360),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(1360),
            data_im_out => mul_im_out(1360)
        );

 
    UMUL_1361 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1361),
            data_im_in => first_stage_im_out(1361),
            re_multiplicator => "0001110101001101", --- 0.457824707031 + j-0.889038085938
            im_multiplicator => "1100011100011010",
            data_re_out => mul_re_out(1361),
            data_im_out => mul_im_out(1361)
        );

 
    UMUL_1362 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1362),
            data_im_in => first_stage_im_out(1362),
            re_multiplicator => "0001100110010011", --- 0.399597167969 + j-0.916687011719
            im_multiplicator => "1100010101010101",
            data_re_out => mul_re_out(1362),
            data_im_out => mul_im_out(1362)
        );

 
    UMUL_1363 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1363),
            data_im_in => first_stage_im_out(1363),
            re_multiplicator => "0001010110111111", --- 0.339782714844 + j-0.940490722656
            im_multiplicator => "1100001111001111",
            data_re_out => mul_re_out(1363),
            data_im_out => mul_im_out(1363)
        );

 
    UMUL_1364 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1364),
            data_im_in => first_stage_im_out(1364),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(1364),
            data_im_out => mul_im_out(1364)
        );

 
    UMUL_1365 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1365),
            data_im_in => first_stage_im_out(1365),
            re_multiplicator => "0000110111010101", --- 0.216125488281 + j-0.976379394531
            im_multiplicator => "1100000110000011",
            data_re_out => mul_re_out(1365),
            data_im_out => mul_im_out(1365)
        );

 
    UMUL_1366 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1366),
            data_im_in => first_stage_im_out(1366),
            re_multiplicator => "0000100111000111", --- 0.152770996094 + j-0.98828125
            im_multiplicator => "1100000011000000",
            data_re_out => mul_re_out(1366),
            data_im_out => mul_im_out(1366)
        );

 
    UMUL_1367 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1367),
            data_im_in => first_stage_im_out(1367),
            re_multiplicator => "0000010110110000", --- 0.0888671875 + j-0.996032714844
            im_multiplicator => "1100000001000001",
            data_re_out => mul_re_out(1367),
            data_im_out => mul_im_out(1367)
        );

 
    UMUL_1368 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1368),
            data_im_in => first_stage_im_out(1368),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(1368),
            data_im_out => mul_im_out(1368)
        );

 
    UMUL_1369 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1369),
            data_im_in => first_stage_im_out(1369),
            re_multiplicator => "1111110101110011", --- -0.0398559570312 + j-0.999206542969
            im_multiplicator => "1100000000001101",
            data_re_out => mul_re_out(1369),
            data_im_out => mul_im_out(1369)
        );

 
    UMUL_1370 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1370),
            data_im_in => first_stage_im_out(1370),
            re_multiplicator => "1111100101010110", --- -0.104125976562 + j-0.994567871094
            im_multiplicator => "1100000001011001",
            data_re_out => mul_re_out(1370),
            data_im_out => mul_im_out(1370)
        );

 
    UMUL_1371 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1371),
            data_im_in => first_stage_im_out(1371),
            re_multiplicator => "1111010101000000", --- -0.16796875 + j-0.985778808594
            im_multiplicator => "1100000011101001",
            data_re_out => mul_re_out(1371),
            data_im_out => mul_im_out(1371)
        );

 
    UMUL_1372 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1372),
            data_im_in => first_stage_im_out(1372),
            re_multiplicator => "1111000100110110", --- -0.231079101562 + j-0.972961425781
            im_multiplicator => "1100000110111011",
            data_re_out => mul_re_out(1372),
            data_im_out => mul_im_out(1372)
        );

 
    UMUL_1373 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1373),
            data_im_in => first_stage_im_out(1373),
            re_multiplicator => "1110110100111100", --- -0.293212890625 + j-0.9560546875
            im_multiplicator => "1100001011010000",
            data_re_out => mul_re_out(1373),
            data_im_out => mul_im_out(1373)
        );

 
    UMUL_1374 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1374),
            data_im_in => first_stage_im_out(1374),
            re_multiplicator => "1110100101010101", --- -0.354187011719 + j-0.935180664062
            im_multiplicator => "1100010000100110",
            data_re_out => mul_re_out(1374),
            data_im_out => mul_im_out(1374)
        );

 
    UMUL_1375 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1375),
            data_im_in => first_stage_im_out(1375),
            re_multiplicator => "1110010110000111", --- -0.413635253906 + j-0.910461425781
            im_multiplicator => "1100010110111011",
            data_re_out => mul_re_out(1375),
            data_im_out => mul_im_out(1375)
        );

 
    UMUL_1376 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1376),
            data_im_in => first_stage_im_out(1376),
            re_multiplicator => "1110000111010101", --- -0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(1376),
            data_im_out => mul_im_out(1376)
        );

 
    UMUL_1377 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1377),
            data_im_in => first_stage_im_out(1377),
            re_multiplicator => "1101111001000010", --- -0.527221679688 + j-0.849731445312
            im_multiplicator => "1100100110011110",
            data_re_out => mul_re_out(1377),
            data_im_out => mul_im_out(1377)
        );

 
    UMUL_1378 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1378),
            data_im_in => first_stage_im_out(1378),
            re_multiplicator => "1101101011010100", --- -0.580810546875 + j-0.814025878906
            im_multiplicator => "1100101111100111",
            data_re_out => mul_re_out(1378),
            data_im_out => mul_im_out(1378)
        );

 
    UMUL_1379 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1379),
            data_im_in => first_stage_im_out(1379),
            re_multiplicator => "1101011110001101", --- -0.632019042969 + j-0.774963378906
            im_multiplicator => "1100111001100111",
            data_re_out => mul_re_out(1379),
            data_im_out => mul_im_out(1379)
        );

 
    UMUL_1380 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1380),
            data_im_in => first_stage_im_out(1380),
            re_multiplicator => "1101010001110001", --- -0.680603027344 + j-0.732666015625
            im_multiplicator => "1101000100011100",
            data_re_out => mul_re_out(1380),
            data_im_out => mul_im_out(1380)
        );

 
    UMUL_1381 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1381),
            data_im_in => first_stage_im_out(1381),
            re_multiplicator => "1101000110000011", --- -0.726379394531 + j-0.687316894531
            im_multiplicator => "1101010000000011",
            data_re_out => mul_re_out(1381),
            data_im_out => mul_im_out(1381)
        );

 
    UMUL_1382 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1382),
            data_im_in => first_stage_im_out(1382),
            re_multiplicator => "1100111011000111", --- -0.769104003906 + j-0.639099121094
            im_multiplicator => "1101011100011001",
            data_re_out => mul_re_out(1382),
            data_im_out => mul_im_out(1382)
        );

 
    UMUL_1383 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1383),
            data_im_in => first_stage_im_out(1383),
            re_multiplicator => "1100110000111111", --- -0.808654785156 + j-0.588256835938
            im_multiplicator => "1101101001011010",
            data_re_out => mul_re_out(1383),
            data_im_out => mul_im_out(1383)
        );

 
    UMUL_1384 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1384),
            data_im_in => first_stage_im_out(1384),
            re_multiplicator => "1100100111101110", --- -0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(1384),
            data_im_out => mul_im_out(1384)
        );

 
    UMUL_1385 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1385),
            data_im_in => first_stage_im_out(1385),
            re_multiplicator => "1100011111010110", --- -0.877563476562 + j-0.4794921875
            im_multiplicator => "1110000101010000",
            data_re_out => mul_re_out(1385),
            data_im_out => mul_im_out(1385)
        );

 
    UMUL_1386 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1386),
            data_im_in => first_stage_im_out(1386),
            re_multiplicator => "1100010111111010", --- -0.906616210938 + j-0.421997070312
            im_multiplicator => "1110010011111110",
            data_re_out => mul_re_out(1386),
            data_im_out => mul_im_out(1386)
        );

 
    UMUL_1387 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1387),
            data_im_in => first_stage_im_out(1387),
            re_multiplicator => "1100010001011100", --- -0.931884765625 + j-0.362731933594
            im_multiplicator => "1110100011001001",
            data_re_out => mul_re_out(1387),
            data_im_out => mul_im_out(1387)
        );

 
    UMUL_1388 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1388),
            data_im_in => first_stage_im_out(1388),
            re_multiplicator => "1100001011111101", --- -0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(1388),
            data_im_out => mul_im_out(1388)
        );

 
    UMUL_1389 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1389),
            data_im_in => first_stage_im_out(1389),
            re_multiplicator => "1100000111011111", --- -0.970764160156 + j-0.239990234375
            im_multiplicator => "1111000010100100",
            data_re_out => mul_re_out(1389),
            data_im_out => mul_im_out(1389)
        );

 
    UMUL_1390 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1390),
            data_im_in => first_stage_im_out(1390),
            re_multiplicator => "1100000100000011", --- -0.984191894531 + j-0.177001953125
            im_multiplicator => "1111010010101100",
            data_re_out => mul_re_out(1390),
            data_im_out => mul_im_out(1390)
        );

 
    UMUL_1391 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1391),
            data_im_in => first_stage_im_out(1391),
            re_multiplicator => "1100000001101001", --- -0.993591308594 + j-0.11328125
            im_multiplicator => "1111100011000000",
            data_re_out => mul_re_out(1391),
            data_im_out => mul_im_out(1391)
        );

 
    UMUL_1392 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1392),
            data_im_in => first_stage_im_out(1392),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(1392),
            data_im_out => mul_im_out(1392)
        );

 
    UMUL_1393 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1393),
            data_im_in => first_stage_im_out(1393),
            re_multiplicator => "1100000000000010", --- -0.999877929688 + j0.0153198242188
            im_multiplicator => "0000000011111011",
            data_re_out => mul_re_out(1393),
            data_im_out => mul_im_out(1393)
        );

 
    UMUL_1394 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1394),
            data_im_in => first_stage_im_out(1394),
            re_multiplicator => "1100000000110100", --- -0.996826171875 + j0.0797119140625
            im_multiplicator => "0000010100011010",
            data_re_out => mul_re_out(1394),
            data_im_out => mul_im_out(1394)
        );

 
    UMUL_1395 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1395),
            data_im_in => first_stage_im_out(1395),
            re_multiplicator => "1100000010101010", --- -0.989624023438 + j0.143676757812
            im_multiplicator => "0000100100110010",
            data_re_out => mul_re_out(1395),
            data_im_out => mul_im_out(1395)
        );

 
    UMUL_1396 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1396),
            data_im_in => first_stage_im_out(1396),
            re_multiplicator => "1100000101100011", --- -0.978332519531 + j0.207092285156
            im_multiplicator => "0000110101000001",
            data_re_out => mul_re_out(1396),
            data_im_out => mul_im_out(1396)
        );

 
    UMUL_1397 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1397),
            data_im_in => first_stage_im_out(1397),
            re_multiplicator => "1100001001011111", --- -0.962951660156 + j0.269653320312
            im_multiplicator => "0001000101000010",
            data_re_out => mul_re_out(1397),
            data_im_out => mul_im_out(1397)
        );

 
    UMUL_1398 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1398),
            data_im_in => first_stage_im_out(1398),
            re_multiplicator => "1100001110011100", --- -0.943603515625 + j0.331115722656
            im_multiplicator => "0001010100110001",
            data_re_out => mul_re_out(1398),
            data_im_out => mul_im_out(1398)
        );

 
    UMUL_1399 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1399),
            data_im_in => first_stage_im_out(1399),
            re_multiplicator => "1100010100011010", --- -0.920288085938 + j0.391174316406
            im_multiplicator => "0001100100001001",
            data_re_out => mul_re_out(1399),
            data_im_out => mul_im_out(1399)
        );

 
    UMUL_1400 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1400),
            data_im_in => first_stage_im_out(1400),
            re_multiplicator => "1100011011010101", --- -0.893249511719 + j0.449584960938
            im_multiplicator => "0001110011000110",
            data_re_out => mul_re_out(1400),
            data_im_out => mul_im_out(1400)
        );

 
    UMUL_1401 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1401),
            data_im_in => first_stage_im_out(1401),
            re_multiplicator => "1100100011001110", --- -0.862426757812 + j0.506164550781
            im_multiplicator => "0010000001100101",
            data_re_out => mul_re_out(1401),
            data_im_out => mul_im_out(1401)
        );

 
    UMUL_1402 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1402),
            data_im_in => first_stage_im_out(1402),
            re_multiplicator => "1100101100000001", --- -0.828063964844 + j0.560668945312
            im_multiplicator => "0010001111100010",
            data_re_out => mul_re_out(1402),
            data_im_out => mul_im_out(1402)
        );

 
    UMUL_1403 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1403),
            data_im_in => first_stage_im_out(1403),
            re_multiplicator => "1100110101101101", --- -0.790222167969 + j0.61279296875
            im_multiplicator => "0010011100111000",
            data_re_out => mul_re_out(1403),
            data_im_out => mul_im_out(1403)
        );

 
    UMUL_1404 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1404),
            data_im_in => first_stage_im_out(1404),
            re_multiplicator => "1101000000001110", --- -0.749145507812 + j0.662414550781
            im_multiplicator => "0010101001100101",
            data_re_out => mul_re_out(1404),
            data_im_out => mul_im_out(1404)
        );

 
    UMUL_1405 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1405),
            data_im_in => first_stage_im_out(1405),
            re_multiplicator => "1101001011100010", --- -0.704956054688 + j0.709289550781
            im_multiplicator => "0010110101100101",
            data_re_out => mul_re_out(1405),
            data_im_out => mul_im_out(1405)
        );

 
    UMUL_1406 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1406),
            data_im_in => first_stage_im_out(1406),
            re_multiplicator => "1101010111100110", --- -0.657836914062 + j0.753173828125
            im_multiplicator => "0011000000110100",
            data_re_out => mul_re_out(1406),
            data_im_out => mul_im_out(1406)
        );

 
    UMUL_1407 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1407),
            data_im_in => first_stage_im_out(1407),
            re_multiplicator => "1101100100010111", --- -0.607971191406 + j0.7939453125
            im_multiplicator => "0011001011010000",
            data_re_out => mul_re_out(1407),
            data_im_out => mul_im_out(1407)
        );

 
    UMUL_1408 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1408),
            data_im_in => first_stage_im_out(1408),
            data_re_out => mul_re_out(1408),
            data_im_out => mul_im_out(1408)
        );

 
    UMUL_1409 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1409),
            data_im_in => first_stage_im_out(1409),
            re_multiplicator => "0011111111011011", --- 0.997741699219 + j-0.0674438476562
            im_multiplicator => "1111101110101111",
            data_re_out => mul_re_out(1409),
            data_im_out => mul_im_out(1409)
        );

 
    UMUL_1410 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1410),
            data_im_in => first_stage_im_out(1410),
            re_multiplicator => "0011111101101011", --- 0.990905761719 + j-0.134582519531
            im_multiplicator => "1111011101100011",
            data_re_out => mul_re_out(1410),
            data_im_out => mul_im_out(1410)
        );

 
    UMUL_1411 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1411),
            data_im_in => first_stage_im_out(1411),
            re_multiplicator => "0011111010110001", --- 0.979553222656 + j-0.201110839844
            im_multiplicator => "1111001100100001",
            data_re_out => mul_re_out(1411),
            data_im_out => mul_im_out(1411)
        );

 
    UMUL_1412 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1412),
            data_im_in => first_stage_im_out(1412),
            re_multiplicator => "0011110110101111", --- 0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(1412),
            data_im_out => mul_im_out(1412)
        );

 
    UMUL_1413 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1413),
            data_im_in => first_stage_im_out(1413),
            re_multiplicator => "0011110001100100", --- 0.943603515625 + j-0.331115722656
            im_multiplicator => "1110101011001111",
            data_re_out => mul_re_out(1413),
            data_im_out => mul_im_out(1413)
        );

 
    UMUL_1414 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1414),
            data_im_in => first_stage_im_out(1414),
            re_multiplicator => "0011101011010011", --- 0.919128417969 + j-0.393981933594
            im_multiplicator => "1110011011001001",
            data_re_out => mul_re_out(1414),
            data_im_out => mul_im_out(1414)
        );

 
    UMUL_1415 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1415),
            data_im_in => first_stage_im_out(1415),
            re_multiplicator => "0011100011111101", --- 0.890441894531 + j-0.455078125
            im_multiplicator => "1110001011100000",
            data_re_out => mul_re_out(1415),
            data_im_out => mul_im_out(1415)
        );

 
    UMUL_1416 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1416),
            data_im_in => first_stage_im_out(1416),
            re_multiplicator => "0011011011100101", --- 0.857727050781 + j-0.514099121094
            im_multiplicator => "1101111100011001",
            data_re_out => mul_re_out(1416),
            data_im_out => mul_im_out(1416)
        );

 
    UMUL_1417 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1417),
            data_im_in => first_stage_im_out(1417),
            re_multiplicator => "0011010010001101", --- 0.821105957031 + j-0.57080078125
            im_multiplicator => "1101101101111000",
            data_re_out => mul_re_out(1417),
            data_im_out => mul_im_out(1417)
        );

 
    UMUL_1418 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1418),
            data_im_in => first_stage_im_out(1418),
            re_multiplicator => "0011000111111000", --- 0.78076171875 + j-0.624877929688
            im_multiplicator => "1101100000000010",
            data_re_out => mul_re_out(1418),
            data_im_out => mul_im_out(1418)
        );

 
    UMUL_1419 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1419),
            data_im_in => first_stage_im_out(1419),
            re_multiplicator => "0010111100101000", --- 0.73681640625 + j-0.676086425781
            im_multiplicator => "1101010010111011",
            data_re_out => mul_re_out(1419),
            data_im_out => mul_im_out(1419)
        );

 
    UMUL_1420 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1420),
            data_im_in => first_stage_im_out(1420),
            re_multiplicator => "0010110000100001", --- 0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(1420),
            data_im_out => mul_im_out(1420)
        );

 
    UMUL_1421 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1421),
            data_im_in => first_stage_im_out(1421),
            re_multiplicator => "0010100011100111", --- 0.639099121094 + j-0.769104003906
            im_multiplicator => "1100111011000111",
            data_re_out => mul_re_out(1421),
            data_im_out => mul_im_out(1421)
        );

 
    UMUL_1422 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1422),
            data_im_in => first_stage_im_out(1422),
            re_multiplicator => "0010010101111110", --- 0.585815429688 + j-0.810485839844
            im_multiplicator => "1100110000100001",
            data_re_out => mul_re_out(1422),
            data_im_out => mul_im_out(1422)
        );

 
    UMUL_1423 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1423),
            data_im_in => first_stage_im_out(1423),
            re_multiplicator => "0010000111101000", --- 0.52978515625 + j-0.84814453125
            im_multiplicator => "1100100110111000",
            data_re_out => mul_re_out(1423),
            data_im_out => mul_im_out(1423)
        );

 
    UMUL_1424 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1424),
            data_im_in => first_stage_im_out(1424),
            re_multiplicator => "0001111000101011", --- 0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(1424),
            data_im_out => mul_im_out(1424)
        );

 
    UMUL_1425 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1425),
            data_im_in => first_stage_im_out(1425),
            re_multiplicator => "0001101001001011", --- 0.410827636719 + j-0.911682128906
            im_multiplicator => "1100010110100111",
            data_re_out => mul_re_out(1425),
            data_im_out => mul_im_out(1425)
        );

 
    UMUL_1426 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1426),
            data_im_in => first_stage_im_out(1426),
            re_multiplicator => "0001011001001100", --- 0.348388671875 + j-0.937316894531
            im_multiplicator => "1100010000000011",
            data_re_out => mul_re_out(1426),
            data_im_out => mul_im_out(1426)
        );

 
    UMUL_1427 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1427),
            data_im_in => first_stage_im_out(1427),
            re_multiplicator => "0001001000110100", --- 0.284423828125 + j-0.958679199219
            im_multiplicator => "1100001010100101",
            data_re_out => mul_re_out(1427),
            data_im_out => mul_im_out(1427)
        );

 
    UMUL_1428 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1428),
            data_im_in => first_stage_im_out(1428),
            re_multiplicator => "0000111000000110", --- 0.219116210938 + j-0.975708007812
            im_multiplicator => "1100000110001110",
            data_re_out => mul_re_out(1428),
            data_im_out => mul_im_out(1428)
        );

 
    UMUL_1429 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1429),
            data_im_in => first_stage_im_out(1429),
            re_multiplicator => "0000100111000111", --- 0.152770996094 + j-0.98828125
            im_multiplicator => "1100000011000000",
            data_re_out => mul_re_out(1429),
            data_im_out => mul_im_out(1429)
        );

 
    UMUL_1430 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1430),
            data_im_in => first_stage_im_out(1430),
            re_multiplicator => "0000010101111110", --- 0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(1430),
            data_im_out => mul_im_out(1430)
        );

 
    UMUL_1431 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1431),
            data_im_in => first_stage_im_out(1431),
            re_multiplicator => "0000000100101110", --- 0.0184326171875 + j-0.999816894531
            im_multiplicator => "1100000000000011",
            data_re_out => mul_re_out(1431),
            data_im_out => mul_im_out(1431)
        );

 
    UMUL_1432 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1432),
            data_im_in => first_stage_im_out(1432),
            re_multiplicator => "1111110011011100", --- -0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(1432),
            data_im_out => mul_im_out(1432)
        );

 
    UMUL_1433 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1433),
            data_im_in => first_stage_im_out(1433),
            re_multiplicator => "1111100010001110", --- -0.116333007812 + j-0.993225097656
            im_multiplicator => "1100000001101111",
            data_re_out => mul_re_out(1433),
            data_im_out => mul_im_out(1433)
        );

 
    UMUL_1434 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1434),
            data_im_in => first_stage_im_out(1434),
            re_multiplicator => "1111010001001001", --- -0.183044433594 + j-0.983093261719
            im_multiplicator => "1100000100010101",
            data_re_out => mul_re_out(1434),
            data_im_out => mul_im_out(1434)
        );

 
    UMUL_1435 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1435),
            data_im_in => first_stage_im_out(1435),
            re_multiplicator => "1111000000010010", --- -0.248901367188 + j-0.968505859375
            im_multiplicator => "1100001000000100",
            data_re_out => mul_re_out(1435),
            data_im_out => mul_im_out(1435)
        );

 
    UMUL_1436 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1436),
            data_im_in => first_stage_im_out(1436),
            re_multiplicator => "1110101111101101", --- -0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(1436),
            data_im_out => mul_im_out(1436)
        );

 
    UMUL_1437 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1437),
            data_im_in => first_stage_im_out(1437),
            re_multiplicator => "1110011111011111", --- -0.377014160156 + j-0.926208496094
            im_multiplicator => "1100010010111001",
            data_re_out => mul_re_out(1437),
            data_im_out => mul_im_out(1437)
        );

 
    UMUL_1438 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1438),
            data_im_in => first_stage_im_out(1438),
            re_multiplicator => "1110001111101110", --- -0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(1438),
            data_im_out => mul_im_out(1438)
        );

 
    UMUL_1439 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1439),
            data_im_in => first_stage_im_out(1439),
            re_multiplicator => "1110000000011101", --- -0.498229980469 + j-0.867065429688
            im_multiplicator => "1100100010000010",
            data_re_out => mul_re_out(1439),
            data_im_out => mul_im_out(1439)
        );

 
    UMUL_1440 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1440),
            data_im_in => first_stage_im_out(1440),
            re_multiplicator => "1101110001110010", --- -0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(1440),
            data_im_out => mul_im_out(1440)
        );

 
    UMUL_1441 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1441),
            data_im_in => first_stage_im_out(1441),
            re_multiplicator => "1101100011101111", --- -0.610412597656 + j-0.792114257812
            im_multiplicator => "1100110101001110",
            data_re_out => mul_re_out(1441),
            data_im_out => mul_im_out(1441)
        );

 
    UMUL_1442 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1442),
            data_im_in => first_stage_im_out(1442),
            re_multiplicator => "1101010110011011", --- -0.662414550781 + j-0.749145507812
            im_multiplicator => "1101000000001110",
            data_re_out => mul_re_out(1442),
            data_im_out => mul_im_out(1442)
        );

 
    UMUL_1443 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1443),
            data_im_in => first_stage_im_out(1443),
            re_multiplicator => "1101001001111000", --- -0.71142578125 + j-0.702758789062
            im_multiplicator => "1101001100000110",
            data_re_out => mul_re_out(1443),
            data_im_out => mul_im_out(1443)
        );

 
    UMUL_1444 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1444),
            data_im_in => first_stage_im_out(1444),
            re_multiplicator => "1100111110001010", --- -0.757202148438 + j-0.653198242188
            im_multiplicator => "1101011000110010",
            data_re_out => mul_re_out(1444),
            data_im_out => mul_im_out(1444)
        );

 
    UMUL_1445 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1445),
            data_im_in => first_stage_im_out(1445),
            re_multiplicator => "1100110011010100", --- -0.799560546875 + j-0.600646972656
            im_multiplicator => "1101100110001111",
            data_re_out => mul_re_out(1445),
            data_im_out => mul_im_out(1445)
        );

 
    UMUL_1446 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1446),
            data_im_in => first_stage_im_out(1446),
            re_multiplicator => "1100101001011011", --- -0.838195800781 + j-0.545349121094
            im_multiplicator => "1101110100011001",
            data_re_out => mul_re_out(1446),
            data_im_out => mul_im_out(1446)
        );

 
    UMUL_1447 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1447),
            data_im_in => first_stage_im_out(1447),
            re_multiplicator => "1100100000011111", --- -0.873107910156 + j-0.487548828125
            im_multiplicator => "1110000011001100",
            data_re_out => mul_re_out(1447),
            data_im_out => mul_im_out(1447)
        );

 
    UMUL_1448 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1448),
            data_im_in => first_stage_im_out(1448),
            re_multiplicator => "1100011000100101", --- -0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(1448),
            data_im_out => mul_im_out(1448)
        );

 
    UMUL_1449 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1449),
            data_im_in => first_stage_im_out(1449),
            re_multiplicator => "1100010001101110", --- -0.930786132812 + j-0.365600585938
            im_multiplicator => "1110100010011010",
            data_re_out => mul_re_out(1449),
            data_im_out => mul_im_out(1449)
        );

 
    UMUL_1450 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1450),
            data_im_in => first_stage_im_out(1450),
            re_multiplicator => "1100001011111101", --- -0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(1450),
            data_im_out => mul_im_out(1450)
        );

 
    UMUL_1451 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1451),
            data_im_in => first_stage_im_out(1451),
            re_multiplicator => "1100000111010011", --- -0.971496582031 + j-0.236999511719
            im_multiplicator => "1111000011010101",
            data_re_out => mul_re_out(1451),
            data_im_out => mul_im_out(1451)
        );

 
    UMUL_1452 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1452),
            data_im_in => first_stage_im_out(1452),
            re_multiplicator => "1100000011110001", --- -0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(1452),
            data_im_out => mul_im_out(1452)
        );

 
    UMUL_1453 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1453),
            data_im_in => first_stage_im_out(1453),
            re_multiplicator => "1100000001011001", --- -0.994567871094 + j-0.104125976562
            im_multiplicator => "1111100101010110",
            data_re_out => mul_re_out(1453),
            data_im_out => mul_im_out(1453)
        );

 
    UMUL_1454 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1454),
            data_im_in => first_stage_im_out(1454),
            re_multiplicator => "1100000000001011", --- -0.999328613281 + j-0.0368041992188
            im_multiplicator => "1111110110100101",
            data_re_out => mul_re_out(1454),
            data_im_out => mul_im_out(1454)
        );

 
    UMUL_1455 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1455),
            data_im_in => first_stage_im_out(1455),
            re_multiplicator => "1100000000001000", --- -0.99951171875 + j0.0307006835938
            im_multiplicator => "0000000111110111",
            data_re_out => mul_re_out(1455),
            data_im_out => mul_im_out(1455)
        );

 
    UMUL_1456 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1456),
            data_im_in => first_stage_im_out(1456),
            re_multiplicator => "1100000001001111", --- -0.995178222656 + j0.0980224609375
            im_multiplicator => "0000011001000110",
            data_re_out => mul_re_out(1456),
            data_im_out => mul_im_out(1456)
        );

 
    UMUL_1457 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1457),
            data_im_in => first_stage_im_out(1457),
            re_multiplicator => "1100000011100000", --- -0.986328125 + j0.164916992188
            im_multiplicator => "0000101010001110",
            data_re_out => mul_re_out(1457),
            data_im_out => mul_im_out(1457)
        );

 
    UMUL_1458 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1458),
            data_im_in => first_stage_im_out(1458),
            re_multiplicator => "1100000110111011", --- -0.972961425781 + j0.231079101562
            im_multiplicator => "0000111011001010",
            data_re_out => mul_re_out(1458),
            data_im_out => mul_im_out(1458)
        );

 
    UMUL_1459 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1459),
            data_im_in => first_stage_im_out(1459),
            re_multiplicator => "1100001011011111", --- -0.955139160156 + j0.296142578125
            im_multiplicator => "0001001011110100",
            data_re_out => mul_re_out(1459),
            data_im_out => mul_im_out(1459)
        );

 
    UMUL_1460 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1460),
            data_im_in => first_stage_im_out(1460),
            re_multiplicator => "1100010001001010", --- -0.932983398438 + j0.359924316406
            im_multiplicator => "0001011100001001",
            data_re_out => mul_re_out(1460),
            data_im_out => mul_im_out(1460)
        );

 
    UMUL_1461 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1461),
            data_im_in => first_stage_im_out(1461),
            re_multiplicator => "1100010111111010", --- -0.906616210938 + j0.421997070312
            im_multiplicator => "0001101100000010",
            data_re_out => mul_re_out(1461),
            data_im_out => mul_im_out(1461)
        );

 
    UMUL_1462 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1462),
            data_im_in => first_stage_im_out(1462),
            re_multiplicator => "1100011111101110", --- -0.876098632812 + j0.482177734375
            im_multiplicator => "0001111011011100",
            data_re_out => mul_re_out(1462),
            data_im_out => mul_im_out(1462)
        );

 
    UMUL_1463 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1463),
            data_im_in => first_stage_im_out(1463),
            re_multiplicator => "1100101000100100", --- -0.841552734375 + j0.540161132812
            im_multiplicator => "0010001010010010",
            data_re_out => mul_re_out(1463),
            data_im_out => mul_im_out(1463)
        );

 
    UMUL_1464 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1464),
            data_im_in => first_stage_im_out(1464),
            re_multiplicator => "1100110010011000", --- -0.80322265625 + j0.595703125
            im_multiplicator => "0010011000100000",
            data_re_out => mul_re_out(1464),
            data_im_out => mul_im_out(1464)
        );

 
    UMUL_1465 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1465),
            data_im_in => first_stage_im_out(1465),
            re_multiplicator => "1100111101001000", --- -0.76123046875 + j0.648498535156
            im_multiplicator => "0010100110000001",
            data_re_out => mul_re_out(1465),
            data_im_out => mul_im_out(1465)
        );

 
    UMUL_1466 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1466),
            data_im_in => first_stage_im_out(1466),
            re_multiplicator => "1101001000110001", --- -0.715759277344 + j0.698364257812
            im_multiplicator => "0010110010110010",
            data_re_out => mul_re_out(1466),
            data_im_out => mul_im_out(1466)
        );

 
    UMUL_1467 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1467),
            data_im_in => first_stage_im_out(1467),
            re_multiplicator => "1101010101010000", --- -0.6669921875 + j0.745056152344
            im_multiplicator => "0010111110101111",
            data_re_out => mul_re_out(1467),
            data_im_out => mul_im_out(1467)
        );

 
    UMUL_1468 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1468),
            data_im_in => first_stage_im_out(1468),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j0.788330078125
            im_multiplicator => "0011001001110100",
            data_re_out => mul_re_out(1468),
            data_im_out => mul_im_out(1468)
        );

 
    UMUL_1469 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1469),
            data_im_in => first_stage_im_out(1469),
            re_multiplicator => "1101110000011110", --- -0.560668945312 + j0.828063964844
            im_multiplicator => "0011010011111111",
            data_re_out => mul_re_out(1469),
            data_im_out => mul_im_out(1469)
        );

 
    UMUL_1470 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1470),
            data_im_in => first_stage_im_out(1470),
            re_multiplicator => "1101111111000110", --- -0.503540039062 + j0.863952636719
            im_multiplicator => "0011011101001011",
            data_re_out => mul_re_out(1470),
            data_im_out => mul_im_out(1470)
        );

 
    UMUL_1471 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1471),
            data_im_in => first_stage_im_out(1471),
            re_multiplicator => "1110001110010100", --- -0.444091796875 + j0.89599609375
            im_multiplicator => "0011100101011000",
            data_re_out => mul_re_out(1471),
            data_im_out => mul_im_out(1471)
        );

 
    UMUL_1472 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1472),
            data_im_in => first_stage_im_out(1472),
            data_re_out => mul_re_out(1472),
            data_im_out => mul_im_out(1472)
        );

 
    UMUL_1473 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1473),
            data_im_in => first_stage_im_out(1473),
            re_multiplicator => "0011111111010111", --- 0.997497558594 + j-0.0704956054688
            im_multiplicator => "1111101101111101",
            data_re_out => mul_re_out(1473),
            data_im_out => mul_im_out(1473)
        );

 
    UMUL_1474 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1474),
            data_im_in => first_stage_im_out(1474),
            re_multiplicator => "0011111101011101", --- 0.990051269531 + j-0.140686035156
            im_multiplicator => "1111011011111111",
            data_re_out => mul_re_out(1474),
            data_im_out => mul_im_out(1474)
        );

 
    UMUL_1475 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1475),
            data_im_in => first_stage_im_out(1475),
            re_multiplicator => "0011111010010010", --- 0.977661132812 + j-0.210083007812
            im_multiplicator => "1111001010001110",
            data_re_out => mul_re_out(1475),
            data_im_out => mul_im_out(1475)
        );

 
    UMUL_1476 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1476),
            data_im_in => first_stage_im_out(1476),
            re_multiplicator => "0011110101111000", --- 0.96044921875 + j-0.278503417969
            im_multiplicator => "1110111000101101",
            data_re_out => mul_re_out(1476),
            data_im_out => mul_im_out(1476)
        );

 
    UMUL_1477 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1477),
            data_im_in => first_stage_im_out(1477),
            re_multiplicator => "0011110000001111", --- 0.938415527344 + j-0.345520019531
            im_multiplicator => "1110100111100011",
            data_re_out => mul_re_out(1477),
            data_im_out => mul_im_out(1477)
        );

 
    UMUL_1478 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1478),
            data_im_in => first_stage_im_out(1478),
            re_multiplicator => "0011101001011001", --- 0.911682128906 + j-0.410827636719
            im_multiplicator => "1110010110110101",
            data_re_out => mul_re_out(1478),
            data_im_out => mul_im_out(1478)
        );

 
    UMUL_1479 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1479),
            data_im_in => first_stage_im_out(1479),
            re_multiplicator => "0011100001011010", --- 0.880493164062 + j-0.47412109375
            im_multiplicator => "1110000110101000",
            data_re_out => mul_re_out(1479),
            data_im_out => mul_im_out(1479)
        );

 
    UMUL_1480 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1480),
            data_im_in => first_stage_im_out(1480),
            re_multiplicator => "0011011000010010", --- 0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(1480),
            data_im_out => mul_im_out(1480)
        );

 
    UMUL_1481 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1481),
            data_im_in => first_stage_im_out(1481),
            re_multiplicator => "0011001110000110", --- 0.805053710938 + j-0.59326171875
            im_multiplicator => "1101101000001000",
            data_re_out => mul_re_out(1481),
            data_im_out => mul_im_out(1481)
        );

 
    UMUL_1482 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1482),
            data_im_in => first_stage_im_out(1482),
            re_multiplicator => "0011000010111000", --- 0.76123046875 + j-0.648498535156
            im_multiplicator => "1101011001111111",
            data_re_out => mul_re_out(1482),
            data_im_out => mul_im_out(1482)
        );

 
    UMUL_1483 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1483),
            data_im_in => first_stage_im_out(1483),
            re_multiplicator => "0010110110101011", --- 0.713562011719 + j-0.700561523438
            im_multiplicator => "1101001100101010",
            data_re_out => mul_re_out(1483),
            data_im_out => mul_im_out(1483)
        );

 
    UMUL_1484 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1484),
            data_im_in => first_stage_im_out(1484),
            re_multiplicator => "0010101001100101", --- 0.662414550781 + j-0.749145507812
            im_multiplicator => "1101000000001110",
            data_re_out => mul_re_out(1484),
            data_im_out => mul_im_out(1484)
        );

 
    UMUL_1485 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1485),
            data_im_in => first_stage_im_out(1485),
            re_multiplicator => "0010011011101001", --- 0.607971191406 + j-0.7939453125
            im_multiplicator => "1100110100110000",
            data_re_out => mul_re_out(1485),
            data_im_out => mul_im_out(1485)
        );

 
    UMUL_1486 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1486),
            data_im_in => first_stage_im_out(1486),
            re_multiplicator => "0010001100111011", --- 0.550476074219 + j-0.834838867188
            im_multiplicator => "1100101010010010",
            data_re_out => mul_re_out(1486),
            data_im_out => mul_im_out(1486)
        );

 
    UMUL_1487 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1487),
            data_im_in => first_stage_im_out(1487),
            re_multiplicator => "0001111101100000", --- 0.490234375 + j-0.87158203125
            im_multiplicator => "1100100000111000",
            data_re_out => mul_re_out(1487),
            data_im_out => mul_im_out(1487)
        );

 
    UMUL_1488 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1488),
            data_im_in => first_stage_im_out(1488),
            re_multiplicator => "0001101101011101", --- 0.427551269531 + j-0.903991699219
            im_multiplicator => "1100011000100101",
            data_re_out => mul_re_out(1488),
            data_im_out => mul_im_out(1488)
        );

 
    UMUL_1489 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1489),
            data_im_in => first_stage_im_out(1489),
            re_multiplicator => "0001011100110111", --- 0.362731933594 + j-0.931884765625
            im_multiplicator => "1100010001011100",
            data_re_out => mul_re_out(1489),
            data_im_out => mul_im_out(1489)
        );

 
    UMUL_1490 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1490),
            data_im_in => first_stage_im_out(1490),
            re_multiplicator => "0001001011110100", --- 0.296142578125 + j-0.955139160156
            im_multiplicator => "1100001011011111",
            data_re_out => mul_re_out(1490),
            data_im_out => mul_im_out(1490)
        );

 
    UMUL_1491 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1491),
            data_im_in => first_stage_im_out(1491),
            re_multiplicator => "0000111010011001", --- 0.228088378906 + j-0.9736328125
            im_multiplicator => "1100000110110000",
            data_re_out => mul_re_out(1491),
            data_im_out => mul_im_out(1491)
        );

 
    UMUL_1492 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1492),
            data_im_in => first_stage_im_out(1492),
            re_multiplicator => "0000101000101011", --- 0.158874511719 + j-0.9873046875
            im_multiplicator => "1100000011010000",
            data_re_out => mul_re_out(1492),
            data_im_out => mul_im_out(1492)
        );

 
    UMUL_1493 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1493),
            data_im_in => first_stage_im_out(1493),
            re_multiplicator => "0000010110110000", --- 0.0888671875 + j-0.996032714844
            im_multiplicator => "1100000001000001",
            data_re_out => mul_re_out(1493),
            data_im_out => mul_im_out(1493)
        );

 
    UMUL_1494 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1494),
            data_im_in => first_stage_im_out(1494),
            re_multiplicator => "0000000100101110", --- 0.0184326171875 + j-0.999816894531
            im_multiplicator => "1100000000000011",
            data_re_out => mul_re_out(1494),
            data_im_out => mul_im_out(1494)
        );

 
    UMUL_1495 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1495),
            data_im_in => first_stage_im_out(1495),
            re_multiplicator => "1111110010101010", --- -0.0521240234375 + j-0.998657226562
            im_multiplicator => "1100000000010110",
            data_re_out => mul_re_out(1495),
            data_im_out => mul_im_out(1495)
        );

 
    UMUL_1496 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1496),
            data_im_in => first_stage_im_out(1496),
            re_multiplicator => "1111100000101010", --- -0.122436523438 + j-0.992492675781
            im_multiplicator => "1100000001111011",
            data_re_out => mul_re_out(1496),
            data_im_out => mul_im_out(1496)
        );

 
    UMUL_1497 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1497),
            data_im_in => first_stage_im_out(1497),
            re_multiplicator => "1111001110110101", --- -0.192077636719 + j-0.981384277344
            im_multiplicator => "1100000100110001",
            data_re_out => mul_re_out(1497),
            data_im_out => mul_im_out(1497)
        );

 
    UMUL_1498 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1498),
            data_im_in => first_stage_im_out(1498),
            re_multiplicator => "1110111101001111", --- -0.260803222656 + j-0.965393066406
            im_multiplicator => "1100001000110111",
            data_re_out => mul_re_out(1498),
            data_im_out => mul_im_out(1498)
        );

 
    UMUL_1499 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1499),
            data_im_in => first_stage_im_out(1499),
            re_multiplicator => "1110101011111111", --- -0.328186035156 + j-0.944580078125
            im_multiplicator => "1100001110001100",
            data_re_out => mul_re_out(1499),
            data_im_out => mul_im_out(1499)
        );

 
    UMUL_1500 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1500),
            data_im_in => first_stage_im_out(1500),
            re_multiplicator => "1110011011001001", --- -0.393981933594 + j-0.919128417969
            im_multiplicator => "1100010100101101",
            data_re_out => mul_re_out(1500),
            data_im_out => mul_im_out(1500)
        );

 
    UMUL_1501 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1501),
            data_im_in => first_stage_im_out(1501),
            re_multiplicator => "1110001010110011", --- -0.457824707031 + j-0.889038085938
            im_multiplicator => "1100011100011010",
            data_re_out => mul_re_out(1501),
            data_im_out => mul_im_out(1501)
        );

 
    UMUL_1502 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1502),
            data_im_in => first_stage_im_out(1502),
            re_multiplicator => "1101111011000011", --- -0.519348144531 + j-0.854553222656
            im_multiplicator => "1100100101001111",
            data_re_out => mul_re_out(1502),
            data_im_out => mul_im_out(1502)
        );

 
    UMUL_1503 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1503),
            data_im_in => first_stage_im_out(1503),
            re_multiplicator => "1101101011111101", --- -0.578308105469 + j-0.815795898438
            im_multiplicator => "1100101111001010",
            data_re_out => mul_re_out(1503),
            data_im_out => mul_im_out(1503)
        );

 
    UMUL_1504 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1504),
            data_im_in => first_stage_im_out(1504),
            re_multiplicator => "1101011101100110", --- -0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(1504),
            data_im_out => mul_im_out(1504)
        );

 
    UMUL_1505 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1505),
            data_im_in => first_stage_im_out(1505),
            re_multiplicator => "1101010000000011", --- -0.687316894531 + j-0.726379394531
            im_multiplicator => "1101000110000011",
            data_re_out => mul_re_out(1505),
            data_im_out => mul_im_out(1505)
        );

 
    UMUL_1506 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1506),
            data_im_in => first_stage_im_out(1506),
            re_multiplicator => "1101000011011000", --- -0.73681640625 + j-0.676086425781
            im_multiplicator => "1101010010111011",
            data_re_out => mul_re_out(1506),
            data_im_out => mul_im_out(1506)
        );

 
    UMUL_1507 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1507),
            data_im_in => first_stage_im_out(1507),
            re_multiplicator => "1100110111101001", --- -0.782653808594 + j-0.622436523438
            im_multiplicator => "1101100000101010",
            data_re_out => mul_re_out(1507),
            data_im_out => mul_im_out(1507)
        );

 
    UMUL_1508 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1508),
            data_im_in => first_stage_im_out(1508),
            re_multiplicator => "1100101100111010", --- -0.824584960938 + j-0.565734863281
            im_multiplicator => "1101101111001011",
            data_re_out => mul_re_out(1508),
            data_im_out => mul_im_out(1508)
        );

 
    UMUL_1509 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1509),
            data_im_in => first_stage_im_out(1509),
            re_multiplicator => "1100100011001110", --- -0.862426757812 + j-0.506164550781
            im_multiplicator => "1101111110011011",
            data_re_out => mul_re_out(1509),
            data_im_out => mul_im_out(1509)
        );

 
    UMUL_1510 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1510),
            data_im_in => first_stage_im_out(1510),
            re_multiplicator => "1100011010101000", --- -0.89599609375 + j-0.444091796875
            im_multiplicator => "1110001110010100",
            data_re_out => mul_re_out(1510),
            data_im_out => mul_im_out(1510)
        );

 
    UMUL_1511 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1511),
            data_im_in => first_stage_im_out(1511),
            re_multiplicator => "1100010011001100", --- -0.925048828125 + j-0.379821777344
            im_multiplicator => "1110011110110001",
            data_re_out => mul_re_out(1511),
            data_im_out => mul_im_out(1511)
        );

 
    UMUL_1512 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1512),
            data_im_in => first_stage_im_out(1512),
            re_multiplicator => "1100001100111011", --- -0.949523925781 + j-0.313659667969
            im_multiplicator => "1110101111101101",
            data_re_out => mul_re_out(1512),
            data_im_out => mul_im_out(1512)
        );

 
    UMUL_1513 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1513),
            data_im_in => first_stage_im_out(1513),
            re_multiplicator => "1100000111110111", --- -0.969299316406 + j-0.245971679688
            im_multiplicator => "1111000001000010",
            data_re_out => mul_re_out(1513),
            data_im_out => mul_im_out(1513)
        );

 
    UMUL_1514 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1514),
            data_im_in => first_stage_im_out(1514),
            re_multiplicator => "1100000100000011", --- -0.984191894531 + j-0.177001953125
            im_multiplicator => "1111010010101100",
            data_re_out => mul_re_out(1514),
            data_im_out => mul_im_out(1514)
        );

 
    UMUL_1515 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1515),
            data_im_in => first_stage_im_out(1515),
            re_multiplicator => "1100000001011110", --- -0.994262695312 + j-0.107177734375
            im_multiplicator => "1111100100100100",
            data_re_out => mul_re_out(1515),
            data_im_out => mul_im_out(1515)
        );

 
    UMUL_1516 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1516),
            data_im_in => first_stage_im_out(1516),
            re_multiplicator => "1100000000001011", --- -0.999328613281 + j-0.0368041992188
            im_multiplicator => "1111110110100101",
            data_re_out => mul_re_out(1516),
            data_im_out => mul_im_out(1516)
        );

 
    UMUL_1517 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1517),
            data_im_in => first_stage_im_out(1517),
            re_multiplicator => "1100000000001001", --- -0.999450683594 + j0.0337524414062
            im_multiplicator => "0000001000101001",
            data_re_out => mul_re_out(1517),
            data_im_out => mul_im_out(1517)
        );

 
    UMUL_1518 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1518),
            data_im_in => first_stage_im_out(1518),
            re_multiplicator => "1100000001011001", --- -0.994567871094 + j0.104125976562
            im_multiplicator => "0000011010101010",
            data_re_out => mul_re_out(1518),
            data_im_out => mul_im_out(1518)
        );

 
    UMUL_1519 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1519),
            data_im_in => first_stage_im_out(1519),
            re_multiplicator => "1100000011111010", --- -0.984741210938 + j0.174011230469
            im_multiplicator => "0000101100100011",
            data_re_out => mul_re_out(1519),
            data_im_out => mul_im_out(1519)
        );

 
    UMUL_1520 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1520),
            data_im_in => first_stage_im_out(1520),
            re_multiplicator => "1100000111101011", --- -0.970031738281 + j0.242980957031
            im_multiplicator => "0000111110001101",
            data_re_out => mul_re_out(1520),
            data_im_out => mul_im_out(1520)
        );

 
    UMUL_1521 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1521),
            data_im_in => first_stage_im_out(1521),
            re_multiplicator => "1100001100101011", --- -0.950500488281 + j0.310791015625
            im_multiplicator => "0001001111100100",
            data_re_out => mul_re_out(1521),
            data_im_out => mul_im_out(1521)
        );

 
    UMUL_1522 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1522),
            data_im_in => first_stage_im_out(1522),
            re_multiplicator => "1100010010111001", --- -0.926208496094 + j0.377014160156
            im_multiplicator => "0001100000100001",
            data_re_out => mul_re_out(1522),
            data_im_out => mul_im_out(1522)
        );

 
    UMUL_1523 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1523),
            data_im_in => first_stage_im_out(1523),
            re_multiplicator => "1100011010010010", --- -0.897338867188 + j0.441345214844
            im_multiplicator => "0001110000111111",
            data_re_out => mul_re_out(1523),
            data_im_out => mul_im_out(1523)
        );

 
    UMUL_1524 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1524),
            data_im_in => first_stage_im_out(1524),
            re_multiplicator => "1100100010110101", --- -0.863952636719 + j0.503540039062
            im_multiplicator => "0010000000111010",
            data_re_out => mul_re_out(1524),
            data_im_out => mul_im_out(1524)
        );

 
    UMUL_1525 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1525),
            data_im_in => first_stage_im_out(1525),
            re_multiplicator => "1100101100011110", --- -0.826293945312 + j0.563171386719
            im_multiplicator => "0010010000001011",
            data_re_out => mul_re_out(1525),
            data_im_out => mul_im_out(1525)
        );

 
    UMUL_1526 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1526),
            data_im_in => first_stage_im_out(1526),
            re_multiplicator => "1100110111001010", --- -0.784545898438 + j0.620056152344
            im_multiplicator => "0010011110101111",
            data_re_out => mul_re_out(1526),
            data_im_out => mul_im_out(1526)
        );

 
    UMUL_1527 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1527),
            data_im_in => first_stage_im_out(1527),
            re_multiplicator => "1101000010110110", --- -0.738891601562 + j0.673828125
            im_multiplicator => "0010101100100000",
            data_re_out => mul_re_out(1527),
            data_im_out => mul_im_out(1527)
        );

 
    UMUL_1528 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1528),
            data_im_in => first_stage_im_out(1528),
            re_multiplicator => "1101001111011111", --- -0.689514160156 + j0.724243164062
            im_multiplicator => "0010111001011010",
            data_re_out => mul_re_out(1528),
            data_im_out => mul_im_out(1528)
        );

 
    UMUL_1529 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1529),
            data_im_in => first_stage_im_out(1529),
            re_multiplicator => "1101011100111111", --- -0.636779785156 + j0.771057128906
            im_multiplicator => "0011000101011001",
            data_re_out => mul_re_out(1529),
            data_im_out => mul_im_out(1529)
        );

 
    UMUL_1530 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1530),
            data_im_in => first_stage_im_out(1530),
            re_multiplicator => "1101101011010100", --- -0.580810546875 + j0.814025878906
            im_multiplicator => "0011010000011001",
            data_re_out => mul_re_out(1530),
            data_im_out => mul_im_out(1530)
        );

 
    UMUL_1531 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1531),
            data_im_in => first_stage_im_out(1531),
            re_multiplicator => "1101111010011000", --- -0.52197265625 + j0.852966308594
            im_multiplicator => "0011011010010111",
            data_re_out => mul_re_out(1531),
            data_im_out => mul_im_out(1531)
        );

 
    UMUL_1532 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1532),
            data_im_in => first_stage_im_out(1532),
            re_multiplicator => "1110001010000111", --- -0.460510253906 + j0.887634277344
            im_multiplicator => "0011100011001111",
            data_re_out => mul_re_out(1532),
            data_im_out => mul_im_out(1532)
        );

 
    UMUL_1533 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1533),
            data_im_in => first_stage_im_out(1533),
            re_multiplicator => "1110011010011011", --- -0.396789550781 + j0.917907714844
            im_multiplicator => "0011101010111111",
            data_re_out => mul_re_out(1533),
            data_im_out => mul_im_out(1533)
        );

 
    UMUL_1534 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1534),
            data_im_in => first_stage_im_out(1534),
            re_multiplicator => "1110101011001111", --- -0.331115722656 + j0.943603515625
            im_multiplicator => "0011110001100100",
            data_re_out => mul_re_out(1534),
            data_im_out => mul_im_out(1534)
        );

 
    UMUL_1535 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1535),
            data_im_in => first_stage_im_out(1535),
            re_multiplicator => "1110111100011111", --- -0.263732910156 + j0.964599609375
            im_multiplicator => "0011110110111100",
            data_re_out => mul_re_out(1535),
            data_im_out => mul_im_out(1535)
        );

 
    UMUL_1536 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1536),
            data_im_in => first_stage_im_out(1536),
            data_re_out => mul_re_out(1536),
            data_im_out => mul_im_out(1536)
        );

 
    UMUL_1537 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1537),
            data_im_in => first_stage_im_out(1537),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(1537),
            data_im_out => mul_im_out(1537)
        );

 
    UMUL_1538 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1538),
            data_im_in => first_stage_im_out(1538),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(1538),
            data_im_out => mul_im_out(1538)
        );

 
    UMUL_1539 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1539),
            data_im_in => first_stage_im_out(1539),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(1539),
            data_im_out => mul_im_out(1539)
        );

 
    UMUL_1540 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1540),
            data_im_in => first_stage_im_out(1540),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(1540),
            data_im_out => mul_im_out(1540)
        );

 
    UMUL_1541 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1541),
            data_im_in => first_stage_im_out(1541),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(1541),
            data_im_out => mul_im_out(1541)
        );

 
    UMUL_1542 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1542),
            data_im_in => first_stage_im_out(1542),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(1542),
            data_im_out => mul_im_out(1542)
        );

 
    UMUL_1543 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1543),
            data_im_in => first_stage_im_out(1543),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(1543),
            data_im_out => mul_im_out(1543)
        );

 
    UMUL_1544 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1544),
            data_im_in => first_stage_im_out(1544),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(1544),
            data_im_out => mul_im_out(1544)
        );

 
    UMUL_1545 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1545),
            data_im_in => first_stage_im_out(1545),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(1545),
            data_im_out => mul_im_out(1545)
        );

 
    UMUL_1546 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1546),
            data_im_in => first_stage_im_out(1546),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(1546),
            data_im_out => mul_im_out(1546)
        );

 
    UMUL_1547 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1547),
            data_im_in => first_stage_im_out(1547),
            re_multiplicator => "0010110000100001", --- 0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(1547),
            data_im_out => mul_im_out(1547)
        );

 
    UMUL_1548 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1548),
            data_im_in => first_stage_im_out(1548),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(1548),
            data_im_out => mul_im_out(1548)
        );

 
    UMUL_1549 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1549),
            data_im_in => first_stage_im_out(1549),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j-0.817565917969
            im_multiplicator => "1100101110101101",
            data_re_out => mul_re_out(1549),
            data_im_out => mul_im_out(1549)
        );

 
    UMUL_1550 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1550),
            data_im_in => first_stage_im_out(1550),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(1550),
            data_im_out => mul_im_out(1550)
        );

 
    UMUL_1551 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1551),
            data_im_in => first_stage_im_out(1551),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(1551),
            data_im_out => mul_im_out(1551)
        );

 
    UMUL_1552 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1552),
            data_im_in => first_stage_im_out(1552),
            re_multiplicator => "0001100001111110", --- 0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(1552),
            data_im_out => mul_im_out(1552)
        );

 
    UMUL_1553 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1553),
            data_im_in => first_stage_im_out(1553),
            re_multiplicator => "0001010000010011", --- 0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(1553),
            data_im_out => mul_im_out(1553)
        );

 
    UMUL_1554 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1554),
            data_im_in => first_stage_im_out(1554),
            re_multiplicator => "0000111110001101", --- 0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(1554),
            data_im_out => mul_im_out(1554)
        );

 
    UMUL_1555 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1555),
            data_im_in => first_stage_im_out(1555),
            re_multiplicator => "0000101011110001", --- 0.170959472656 + j-0.985290527344
            im_multiplicator => "1100000011110001",
            data_re_out => mul_re_out(1555),
            data_im_out => mul_im_out(1555)
        );

 
    UMUL_1556 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1556),
            data_im_in => first_stage_im_out(1556),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(1556),
            data_im_out => mul_im_out(1556)
        );

 
    UMUL_1557 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1557),
            data_im_in => first_stage_im_out(1557),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(1557),
            data_im_out => mul_im_out(1557)
        );

 
    UMUL_1558 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1558),
            data_im_in => first_stage_im_out(1558),
            re_multiplicator => "1111110011011100", --- -0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(1558),
            data_im_out => mul_im_out(1558)
        );

 
    UMUL_1559 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1559),
            data_im_in => first_stage_im_out(1559),
            re_multiplicator => "1111100000101010", --- -0.122436523438 + j-0.992492675781
            im_multiplicator => "1100000001111011",
            data_re_out => mul_re_out(1559),
            data_im_out => mul_im_out(1559)
        );

 
    UMUL_1560 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1560),
            data_im_in => first_stage_im_out(1560),
            re_multiplicator => "1111001110000100", --- -0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(1560),
            data_im_out => mul_im_out(1560)
        );

 
    UMUL_1561 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1561),
            data_im_in => first_stage_im_out(1561),
            re_multiplicator => "1110111011101110", --- -0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(1561),
            data_im_out => mul_im_out(1561)
        );

 
    UMUL_1562 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1562),
            data_im_in => first_stage_im_out(1562),
            re_multiplicator => "1110101001110000", --- -0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(1562),
            data_im_out => mul_im_out(1562)
        );

 
    UMUL_1563 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1563),
            data_im_in => first_stage_im_out(1563),
            re_multiplicator => "1110011000010001", --- -0.405212402344 + j-0.914184570312
            im_multiplicator => "1100010101111110",
            data_re_out => mul_re_out(1563),
            data_im_out => mul_im_out(1563)
        );

 
    UMUL_1564 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1564),
            data_im_in => first_stage_im_out(1564),
            re_multiplicator => "1110000111010101", --- -0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(1564),
            data_im_out => mul_im_out(1564)
        );

 
    UMUL_1565 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1565),
            data_im_in => first_stage_im_out(1565),
            re_multiplicator => "1101110111000011", --- -0.534973144531 + j-0.844848632812
            im_multiplicator => "1100100111101110",
            data_re_out => mul_re_out(1565),
            data_im_out => mul_im_out(1565)
        );

 
    UMUL_1566 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1566),
            data_im_in => first_stage_im_out(1566),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(1566),
            data_im_out => mul_im_out(1566)
        );

 
    UMUL_1567 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1567),
            data_im_in => first_stage_im_out(1567),
            re_multiplicator => "1101011000110010", --- -0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(1567),
            data_im_out => mul_im_out(1567)
        );

 
    UMUL_1568 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1568),
            data_im_in => first_stage_im_out(1568),
            re_multiplicator => "1101001010111111", --- -0.707092285156 + j-0.707092285156
            im_multiplicator => "1101001010111111",
            data_re_out => mul_re_out(1568),
            data_im_out => mul_im_out(1568)
        );

 
    UMUL_1569 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1569),
            data_im_in => first_stage_im_out(1569),
            re_multiplicator => "1100111110001010", --- -0.757202148438 + j-0.653198242188
            im_multiplicator => "1101011000110010",
            data_re_out => mul_re_out(1569),
            data_im_out => mul_im_out(1569)
        );

 
    UMUL_1570 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1570),
            data_im_in => first_stage_im_out(1570),
            re_multiplicator => "1100110010011000", --- -0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(1570),
            data_im_out => mul_im_out(1570)
        );

 
    UMUL_1571 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1571),
            data_im_in => first_stage_im_out(1571),
            re_multiplicator => "1100100111101110", --- -0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(1571),
            data_im_out => mul_im_out(1571)
        );

 
    UMUL_1572 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1572),
            data_im_in => first_stage_im_out(1572),
            re_multiplicator => "1100011110001111", --- -0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(1572),
            data_im_out => mul_im_out(1572)
        );

 
    UMUL_1573 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1573),
            data_im_in => first_stage_im_out(1573),
            re_multiplicator => "1100010101111110", --- -0.914184570312 + j-0.405212402344
            im_multiplicator => "1110011000010001",
            data_re_out => mul_re_out(1573),
            data_im_out => mul_im_out(1573)
        );

 
    UMUL_1574 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1574),
            data_im_in => first_stage_im_out(1574),
            re_multiplicator => "1100001110111110", --- -0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(1574),
            data_im_out => mul_im_out(1574)
        );

 
    UMUL_1575 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1575),
            data_im_in => first_stage_im_out(1575),
            re_multiplicator => "1100001001010001", --- -0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(1575),
            data_im_out => mul_im_out(1575)
        );

 
    UMUL_1576 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1576),
            data_im_in => first_stage_im_out(1576),
            re_multiplicator => "1100000100111011", --- -0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(1576),
            data_im_out => mul_im_out(1576)
        );

 
    UMUL_1577 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1577),
            data_im_in => first_stage_im_out(1577),
            re_multiplicator => "1100000001111011", --- -0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(1577),
            data_im_out => mul_im_out(1577)
        );

 
    UMUL_1578 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1578),
            data_im_in => first_stage_im_out(1578),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(1578),
            data_im_out => mul_im_out(1578)
        );

 
    UMUL_1579 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1579),
            data_im_in => first_stage_im_out(1579),
            re_multiplicator => "1100000000000101", --- -0.999694824219 + j0.0245361328125
            im_multiplicator => "0000000110010010",
            data_re_out => mul_re_out(1579),
            data_im_out => mul_im_out(1579)
        );

 
    UMUL_1580 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1580),
            data_im_in => first_stage_im_out(1580),
            re_multiplicator => "1100000001001111", --- -0.995178222656 + j0.0980224609375
            im_multiplicator => "0000011001000110",
            data_re_out => mul_re_out(1580),
            data_im_out => mul_im_out(1580)
        );

 
    UMUL_1581 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1581),
            data_im_in => first_stage_im_out(1581),
            re_multiplicator => "1100000011110001", --- -0.985290527344 + j0.170959472656
            im_multiplicator => "0000101011110001",
            data_re_out => mul_re_out(1581),
            data_im_out => mul_im_out(1581)
        );

 
    UMUL_1582 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1582),
            data_im_in => first_stage_im_out(1582),
            re_multiplicator => "1100000111101011", --- -0.970031738281 + j0.242980957031
            im_multiplicator => "0000111110001101",
            data_re_out => mul_re_out(1582),
            data_im_out => mul_im_out(1582)
        );

 
    UMUL_1583 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1583),
            data_im_in => first_stage_im_out(1583),
            re_multiplicator => "1100001100111011", --- -0.949523925781 + j0.313659667969
            im_multiplicator => "0001010000010011",
            data_re_out => mul_re_out(1583),
            data_im_out => mul_im_out(1583)
        );

 
    UMUL_1584 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1584),
            data_im_in => first_stage_im_out(1584),
            re_multiplicator => "1100010011011111", --- -0.923889160156 + j0.382690429688
            im_multiplicator => "0001100001111110",
            data_re_out => mul_re_out(1584),
            data_im_out => mul_im_out(1584)
        );

 
    UMUL_1585 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1585),
            data_im_in => first_stage_im_out(1585),
            re_multiplicator => "1100011011010101", --- -0.893249511719 + j0.449584960938
            im_multiplicator => "0001110011000110",
            data_re_out => mul_re_out(1585),
            data_im_out => mul_im_out(1585)
        );

 
    UMUL_1586 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1586),
            data_im_in => first_stage_im_out(1586),
            re_multiplicator => "1100100100011011", --- -0.857727050781 + j0.514099121094
            im_multiplicator => "0010000011100111",
            data_re_out => mul_re_out(1586),
            data_im_out => mul_im_out(1586)
        );

 
    UMUL_1587 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1587),
            data_im_in => first_stage_im_out(1587),
            re_multiplicator => "1100101110101101", --- -0.817565917969 + j0.575805664062
            im_multiplicator => "0010010011011010",
            data_re_out => mul_re_out(1587),
            data_im_out => mul_im_out(1587)
        );

 
    UMUL_1588 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1588),
            data_im_in => first_stage_im_out(1588),
            re_multiplicator => "1100111010000111", --- -0.773010253906 + j0.634399414062
            im_multiplicator => "0010100010011010",
            data_re_out => mul_re_out(1588),
            data_im_out => mul_im_out(1588)
        );

 
    UMUL_1589 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1589),
            data_im_in => first_stage_im_out(1589),
            re_multiplicator => "1101000110100110", --- -0.724243164062 + j0.689514160156
            im_multiplicator => "0010110000100001",
            data_re_out => mul_re_out(1589),
            data_im_out => mul_im_out(1589)
        );

 
    UMUL_1590 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1590),
            data_im_in => first_stage_im_out(1590),
            re_multiplicator => "1101010100000101", --- -0.671569824219 + j0.740966796875
            im_multiplicator => "0010111101101100",
            data_re_out => mul_re_out(1590),
            data_im_out => mul_im_out(1590)
        );

 
    UMUL_1591 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1591),
            data_im_in => first_stage_im_out(1591),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j0.788330078125
            im_multiplicator => "0011001001110100",
            data_re_out => mul_re_out(1591),
            data_im_out => mul_im_out(1591)
        );

 
    UMUL_1592 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1592),
            data_im_in => first_stage_im_out(1592),
            re_multiplicator => "1101110001110010", --- -0.555541992188 + j0.831481933594
            im_multiplicator => "0011010100110111",
            data_re_out => mul_re_out(1592),
            data_im_out => mul_im_out(1592)
        );

 
    UMUL_1593 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1593),
            data_im_in => first_stage_im_out(1593),
            re_multiplicator => "1110000001110100", --- -0.492919921875 + j0.8701171875
            im_multiplicator => "0011011110110000",
            data_re_out => mul_re_out(1593),
            data_im_out => mul_im_out(1593)
        );

 
    UMUL_1594 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1594),
            data_im_in => first_stage_im_out(1594),
            re_multiplicator => "1110010010100011", --- -0.427551269531 + j0.903991699219
            im_multiplicator => "0011100111011011",
            data_re_out => mul_re_out(1594),
            data_im_out => mul_im_out(1594)
        );

 
    UMUL_1595 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1595),
            data_im_in => first_stage_im_out(1595),
            re_multiplicator => "1110100011110111", --- -0.359924316406 + j0.932983398438
            im_multiplicator => "0011101110110110",
            data_re_out => mul_re_out(1595),
            data_im_out => mul_im_out(1595)
        );

 
    UMUL_1596 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1596),
            data_im_in => first_stage_im_out(1596),
            re_multiplicator => "1110110101101100", --- -0.290283203125 + j0.956970214844
            im_multiplicator => "0011110100111111",
            data_re_out => mul_re_out(1596),
            data_im_out => mul_im_out(1596)
        );

 
    UMUL_1597 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1597),
            data_im_in => first_stage_im_out(1597),
            re_multiplicator => "1111000111111010", --- -0.219116210938 + j0.975708007812
            im_multiplicator => "0011111001110010",
            data_re_out => mul_re_out(1597),
            data_im_out => mul_im_out(1597)
        );

 
    UMUL_1598 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1598),
            data_im_in => first_stage_im_out(1598),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j0.989196777344
            im_multiplicator => "0011111101001111",
            data_re_out => mul_re_out(1598),
            data_im_out => mul_im_out(1598)
        );

 
    UMUL_1599 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1599),
            data_im_in => first_stage_im_out(1599),
            re_multiplicator => "1111101101001011", --- -0.0735473632812 + j0.997314453125
            im_multiplicator => "0011111111010100",
            data_re_out => mul_re_out(1599),
            data_im_out => mul_im_out(1599)
        );

 
    UMUL_1600 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1600),
            data_im_in => first_stage_im_out(1600),
            data_re_out => mul_re_out(1600),
            data_im_out => mul_im_out(1600)
        );

 
    UMUL_1601 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1601),
            data_im_in => first_stage_im_out(1601),
            re_multiplicator => "0011111111010000", --- 0.9970703125 + j-0.0765991210938
            im_multiplicator => "1111101100011001",
            data_re_out => mul_re_out(1601),
            data_im_out => mul_im_out(1601)
        );

 
    UMUL_1602 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1602),
            data_im_in => first_stage_im_out(1602),
            re_multiplicator => "0011111101000000", --- 0.98828125 + j-0.152770996094
            im_multiplicator => "1111011000111001",
            data_re_out => mul_re_out(1602),
            data_im_out => mul_im_out(1602)
        );

 
    UMUL_1603 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1603),
            data_im_in => first_stage_im_out(1603),
            re_multiplicator => "0011111001010000", --- 0.9736328125 + j-0.228088378906
            im_multiplicator => "1111000101100111",
            data_re_out => mul_re_out(1603),
            data_im_out => mul_im_out(1603)
        );

 
    UMUL_1604 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1604),
            data_im_in => first_stage_im_out(1604),
            re_multiplicator => "0011110100000011", --- 0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(1604),
            data_im_out => mul_im_out(1604)
        );

 
    UMUL_1605 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1605),
            data_im_in => first_stage_im_out(1605),
            re_multiplicator => "0011101101011010", --- 0.927368164062 + j-0.374145507812
            im_multiplicator => "1110100000001110",
            data_re_out => mul_re_out(1605),
            data_im_out => mul_im_out(1605)
        );

 
    UMUL_1606 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1606),
            data_im_in => first_stage_im_out(1606),
            re_multiplicator => "0011100101011000", --- 0.89599609375 + j-0.444091796875
            im_multiplicator => "1110001110010100",
            data_re_out => mul_re_out(1606),
            data_im_out => mul_im_out(1606)
        );

 
    UMUL_1607 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1607),
            data_im_in => first_stage_im_out(1607),
            re_multiplicator => "0011011011111111", --- 0.859313964844 + j-0.511474609375
            im_multiplicator => "1101111101000100",
            data_re_out => mul_re_out(1607),
            data_im_out => mul_im_out(1607)
        );

 
    UMUL_1608 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1608),
            data_im_in => first_stage_im_out(1608),
            re_multiplicator => "0011010001010011", --- 0.817565917969 + j-0.575805664062
            im_multiplicator => "1101101100100110",
            data_re_out => mul_re_out(1608),
            data_im_out => mul_im_out(1608)
        );

 
    UMUL_1609 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1609),
            data_im_in => first_stage_im_out(1609),
            re_multiplicator => "0011000101011001", --- 0.771057128906 + j-0.636779785156
            im_multiplicator => "1101011100111111",
            data_re_out => mul_re_out(1609),
            data_im_out => mul_im_out(1609)
        );

 
    UMUL_1610 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1610),
            data_im_in => first_stage_im_out(1610),
            re_multiplicator => "0010111000010101", --- 0.720031738281 + j-0.693969726562
            im_multiplicator => "1101001110010110",
            data_re_out => mul_re_out(1610),
            data_im_out => mul_im_out(1610)
        );

 
    UMUL_1611 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1611),
            data_im_in => first_stage_im_out(1611),
            re_multiplicator => "0010101010001011", --- 0.664733886719 + j-0.7470703125
            im_multiplicator => "1101000000110000",
            data_re_out => mul_re_out(1611),
            data_im_out => mul_im_out(1611)
        );

 
    UMUL_1612 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1612),
            data_im_in => first_stage_im_out(1612),
            re_multiplicator => "0010011011000001", --- 0.605529785156 + j-0.795837402344
            im_multiplicator => "1100110100010001",
            data_re_out => mul_re_out(1612),
            data_im_out => mul_im_out(1612)
        );

 
    UMUL_1613 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1613),
            data_im_in => first_stage_im_out(1613),
            re_multiplicator => "0010001010111100", --- 0.542724609375 + j-0.839904785156
            im_multiplicator => "1100101000111111",
            data_re_out => mul_re_out(1613),
            data_im_out => mul_im_out(1613)
        );

 
    UMUL_1614 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1614),
            data_im_in => first_stage_im_out(1614),
            re_multiplicator => "0001111010000100", --- 0.476806640625 + j-0.879028320312
            im_multiplicator => "1100011110111110",
            data_re_out => mul_re_out(1614),
            data_im_out => mul_im_out(1614)
        );

 
    UMUL_1615 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1615),
            data_im_in => first_stage_im_out(1615),
            re_multiplicator => "0001101000011101", --- 0.408020019531 + j-0.912963867188
            im_multiplicator => "1100010110010010",
            data_re_out => mul_re_out(1615),
            data_im_out => mul_im_out(1615)
        );

 
    UMUL_1616 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1616),
            data_im_in => first_stage_im_out(1616),
            re_multiplicator => "0001010110010000", --- 0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(1616),
            data_im_out => mul_im_out(1616)
        );

 
    UMUL_1617 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1617),
            data_im_in => first_stage_im_out(1617),
            re_multiplicator => "0001000011100001", --- 0.263732910156 + j-0.964599609375
            im_multiplicator => "1100001001000100",
            data_re_out => mul_re_out(1617),
            data_im_out => mul_im_out(1617)
        );

 
    UMUL_1618 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1618),
            data_im_in => first_stage_im_out(1618),
            re_multiplicator => "0000110000011010", --- 0.189086914062 + j-0.98193359375
            im_multiplicator => "1100000100101000",
            data_re_out => mul_re_out(1618),
            data_im_out => mul_im_out(1618)
        );

 
    UMUL_1619 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1619),
            data_im_in => first_stage_im_out(1619),
            re_multiplicator => "0000011101000000", --- 0.11328125 + j-0.993591308594
            im_multiplicator => "1100000001101001",
            data_re_out => mul_re_out(1619),
            data_im_out => mul_im_out(1619)
        );

 
    UMUL_1620 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1620),
            data_im_in => first_stage_im_out(1620),
            re_multiplicator => "0000001001011011", --- 0.0368041992188 + j-0.999328613281
            im_multiplicator => "1100000000001011",
            data_re_out => mul_re_out(1620),
            data_im_out => mul_im_out(1620)
        );

 
    UMUL_1621 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1621),
            data_im_in => first_stage_im_out(1621),
            re_multiplicator => "1111110101110011", --- -0.0398559570312 + j-0.999206542969
            im_multiplicator => "1100000000001101",
            data_re_out => mul_re_out(1621),
            data_im_out => mul_im_out(1621)
        );

 
    UMUL_1622 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1622),
            data_im_in => first_stage_im_out(1622),
            re_multiplicator => "1111100010001110", --- -0.116333007812 + j-0.993225097656
            im_multiplicator => "1100000001101111",
            data_re_out => mul_re_out(1622),
            data_im_out => mul_im_out(1622)
        );

 
    UMUL_1623 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1623),
            data_im_in => first_stage_im_out(1623),
            re_multiplicator => "1111001110110101", --- -0.192077636719 + j-0.981384277344
            im_multiplicator => "1100000100110001",
            data_re_out => mul_re_out(1623),
            data_im_out => mul_im_out(1623)
        );

 
    UMUL_1624 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1624),
            data_im_in => first_stage_im_out(1624),
            re_multiplicator => "1110111011101110", --- -0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(1624),
            data_im_out => mul_im_out(1624)
        );

 
    UMUL_1625 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1625),
            data_im_in => first_stage_im_out(1625),
            re_multiplicator => "1110101001000001", --- -0.339782714844 + j-0.940490722656
            im_multiplicator => "1100001111001111",
            data_re_out => mul_re_out(1625),
            data_im_out => mul_im_out(1625)
        );

 
    UMUL_1626 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1626),
            data_im_in => first_stage_im_out(1626),
            re_multiplicator => "1110010110110101", --- -0.410827636719 + j-0.911682128906
            im_multiplicator => "1100010110100111",
            data_re_out => mul_re_out(1626),
            data_im_out => mul_im_out(1626)
        );

 
    UMUL_1627 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1627),
            data_im_in => first_stage_im_out(1627),
            re_multiplicator => "1110000101010000", --- -0.4794921875 + j-0.877563476562
            im_multiplicator => "1100011111010110",
            data_re_out => mul_re_out(1627),
            data_im_out => mul_im_out(1627)
        );

 
    UMUL_1628 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1628),
            data_im_in => first_stage_im_out(1628),
            re_multiplicator => "1101110100011001", --- -0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(1628),
            data_im_out => mul_im_out(1628)
        );

 
    UMUL_1629 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1629),
            data_im_in => first_stage_im_out(1629),
            re_multiplicator => "1101100100010111", --- -0.607971191406 + j-0.7939453125
            im_multiplicator => "1100110100110000",
            data_re_out => mul_re_out(1629),
            data_im_out => mul_im_out(1629)
        );

 
    UMUL_1630 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1630),
            data_im_in => first_stage_im_out(1630),
            re_multiplicator => "1101010101010000", --- -0.6669921875 + j-0.745056152344
            im_multiplicator => "1101000001010001",
            data_re_out => mul_re_out(1630),
            data_im_out => mul_im_out(1630)
        );

 
    UMUL_1631 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1631),
            data_im_in => first_stage_im_out(1631),
            re_multiplicator => "1101000111001001", --- -0.722106933594 + j-0.691772460938
            im_multiplicator => "1101001110111010",
            data_re_out => mul_re_out(1631),
            data_im_out => mul_im_out(1631)
        );

 
    UMUL_1632 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1632),
            data_im_in => first_stage_im_out(1632),
            re_multiplicator => "1100111010000111", --- -0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(1632),
            data_im_out => mul_im_out(1632)
        );

 
    UMUL_1633 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1633),
            data_im_in => first_stage_im_out(1633),
            re_multiplicator => "1100101110010000", --- -0.8193359375 + j-0.573303222656
            im_multiplicator => "1101101101001111",
            data_re_out => mul_re_out(1633),
            data_im_out => mul_im_out(1633)
        );

 
    UMUL_1634 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1634),
            data_im_in => first_stage_im_out(1634),
            re_multiplicator => "1100100011101000", --- -0.86083984375 + j-0.508850097656
            im_multiplicator => "1101111101101111",
            data_re_out => mul_re_out(1634),
            data_im_out => mul_im_out(1634)
        );

 
    UMUL_1635 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1635),
            data_im_in => first_stage_im_out(1635),
            re_multiplicator => "1100011010010010", --- -0.897338867188 + j-0.441345214844
            im_multiplicator => "1110001111000001",
            data_re_out => mul_re_out(1635),
            data_im_out => mul_im_out(1635)
        );

 
    UMUL_1636 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1636),
            data_im_in => first_stage_im_out(1636),
            re_multiplicator => "1100010010010011", --- -0.928527832031 + j-0.371337890625
            im_multiplicator => "1110100000111100",
            data_re_out => mul_re_out(1636),
            data_im_out => mul_im_out(1636)
        );

 
    UMUL_1637 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1637),
            data_im_in => first_stage_im_out(1637),
            re_multiplicator => "1100001011101110", --- -0.954223632812 + j-0.299072265625
            im_multiplicator => "1110110011011100",
            data_re_out => mul_re_out(1637),
            data_im_out => mul_im_out(1637)
        );

 
    UMUL_1638 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1638),
            data_im_in => first_stage_im_out(1638),
            re_multiplicator => "1100000110100100", --- -0.974365234375 + j-0.22509765625
            im_multiplicator => "1111000110011000",
            data_re_out => mul_re_out(1638),
            data_im_out => mul_im_out(1638)
        );

 
    UMUL_1639 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1639),
            data_im_in => first_stage_im_out(1639),
            re_multiplicator => "1100000010111001", --- -0.988708496094 + j-0.149780273438
            im_multiplicator => "1111011001101010",
            data_re_out => mul_re_out(1639),
            data_im_out => mul_im_out(1639)
        );

 
    UMUL_1640 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1640),
            data_im_in => first_stage_im_out(1640),
            re_multiplicator => "1100000000101100", --- -0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(1640),
            data_im_out => mul_im_out(1640)
        );

 
    UMUL_1641 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1641),
            data_im_in => first_stage_im_out(1641),
            re_multiplicator => "1100000000000000", --- -1.0 + j0.0030517578125
            im_multiplicator => "0000000000110010",
            data_re_out => mul_re_out(1641),
            data_im_out => mul_im_out(1641)
        );

 
    UMUL_1642 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1642),
            data_im_in => first_stage_im_out(1642),
            re_multiplicator => "1100000000110100", --- -0.996826171875 + j0.0797119140625
            im_multiplicator => "0000010100011010",
            data_re_out => mul_re_out(1642),
            data_im_out => mul_im_out(1642)
        );

 
    UMUL_1643 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1643),
            data_im_in => first_stage_im_out(1643),
            re_multiplicator => "1100000011001000", --- -0.98779296875 + j0.155822753906
            im_multiplicator => "0000100111111001",
            data_re_out => mul_re_out(1643),
            data_im_out => mul_im_out(1643)
        );

 
    UMUL_1644 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1644),
            data_im_in => first_stage_im_out(1644),
            re_multiplicator => "1100000110111011", --- -0.972961425781 + j0.231079101562
            im_multiplicator => "0000111011001010",
            data_re_out => mul_re_out(1644),
            data_im_out => mul_im_out(1644)
        );

 
    UMUL_1645 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1645),
            data_im_in => first_stage_im_out(1645),
            re_multiplicator => "1100001100001100", --- -0.952392578125 + j0.304931640625
            im_multiplicator => "0001001110000100",
            data_re_out => mul_re_out(1645),
            data_im_out => mul_im_out(1645)
        );

 
    UMUL_1646 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1646),
            data_im_in => first_stage_im_out(1646),
            re_multiplicator => "1100010010111001", --- -0.926208496094 + j0.377014160156
            im_multiplicator => "0001100000100001",
            data_re_out => mul_re_out(1646),
            data_im_out => mul_im_out(1646)
        );

 
    UMUL_1647 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1647),
            data_im_in => first_stage_im_out(1647),
            re_multiplicator => "1100011010111111", --- -0.894592285156 + j0.446838378906
            im_multiplicator => "0001110010011001",
            data_re_out => mul_re_out(1647),
            data_im_out => mul_im_out(1647)
        );

 
    UMUL_1648 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1648),
            data_im_in => first_stage_im_out(1648),
            re_multiplicator => "1100100100011011", --- -0.857727050781 + j0.514099121094
            im_multiplicator => "0010000011100111",
            data_re_out => mul_re_out(1648),
            data_im_out => mul_im_out(1648)
        );

 
    UMUL_1649 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1649),
            data_im_in => first_stage_im_out(1649),
            re_multiplicator => "1100101111001010", --- -0.815795898438 + j0.578308105469
            im_multiplicator => "0010010100000011",
            data_re_out => mul_re_out(1649),
            data_im_out => mul_im_out(1649)
        );

 
    UMUL_1650 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1650),
            data_im_in => first_stage_im_out(1650),
            re_multiplicator => "1100111011000111", --- -0.769104003906 + j0.639099121094
            im_multiplicator => "0010100011100111",
            data_re_out => mul_re_out(1650),
            data_im_out => mul_im_out(1650)
        );

 
    UMUL_1651 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1651),
            data_im_in => first_stage_im_out(1651),
            re_multiplicator => "1101001000001110", --- -0.717895507812 + j0.696166992188
            im_multiplicator => "0010110010001110",
            data_re_out => mul_re_out(1651),
            data_im_out => mul_im_out(1651)
        );

 
    UMUL_1652 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1652),
            data_im_in => first_stage_im_out(1652),
            re_multiplicator => "1101010110011011", --- -0.662414550781 + j0.749145507812
            im_multiplicator => "0010111111110010",
            data_re_out => mul_re_out(1652),
            data_im_out => mul_im_out(1652)
        );

 
    UMUL_1653 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1653),
            data_im_in => first_stage_im_out(1653),
            re_multiplicator => "1101100101100111", --- -0.603088378906 + j0.797668457031
            im_multiplicator => "0011001100001101",
            data_re_out => mul_re_out(1653),
            data_im_out => mul_im_out(1653)
        );

 
    UMUL_1654 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1654),
            data_im_in => first_stage_im_out(1654),
            re_multiplicator => "1101110101101110", --- -0.540161132812 + j0.841552734375
            im_multiplicator => "0011010111011100",
            data_re_out => mul_re_out(1654),
            data_im_out => mul_im_out(1654)
        );

 
    UMUL_1655 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1655),
            data_im_in => first_stage_im_out(1655),
            re_multiplicator => "1110000110101000", --- -0.47412109375 + j0.880493164062
            im_multiplicator => "0011100001011010",
            data_re_out => mul_re_out(1655),
            data_im_out => mul_im_out(1655)
        );

 
    UMUL_1656 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1656),
            data_im_in => first_stage_im_out(1656),
            re_multiplicator => "1110011000010001", --- -0.405212402344 + j0.914184570312
            im_multiplicator => "0011101010000010",
            data_re_out => mul_re_out(1656),
            data_im_out => mul_im_out(1656)
        );

 
    UMUL_1657 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1657),
            data_im_in => first_stage_im_out(1657),
            re_multiplicator => "1110101010100000", --- -0.333984375 + j0.942565917969
            im_multiplicator => "0011110001010011",
            data_re_out => mul_re_out(1657),
            data_im_out => mul_im_out(1657)
        );

 
    UMUL_1658 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1658),
            data_im_in => first_stage_im_out(1658),
            re_multiplicator => "1110111101001111", --- -0.260803222656 + j0.965393066406
            im_multiplicator => "0011110111001001",
            data_re_out => mul_re_out(1658),
            data_im_out => mul_im_out(1658)
        );

 
    UMUL_1659 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1659),
            data_im_in => first_stage_im_out(1659),
            re_multiplicator => "1111010000011000", --- -0.18603515625 + j0.982543945312
            im_multiplicator => "0011111011100010",
            data_re_out => mul_re_out(1659),
            data_im_out => mul_im_out(1659)
        );

 
    UMUL_1660 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1660),
            data_im_in => first_stage_im_out(1660),
            re_multiplicator => "1111100011110010", --- -0.110229492188 + j0.993896484375
            im_multiplicator => "0011111110011100",
            data_re_out => mul_re_out(1660),
            data_im_out => mul_im_out(1660)
        );

 
    UMUL_1661 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1661),
            data_im_in => first_stage_im_out(1661),
            re_multiplicator => "1111110111010111", --- -0.0337524414062 + j0.999450683594
            im_multiplicator => "0011111111110111",
            data_re_out => mul_re_out(1661),
            data_im_out => mul_im_out(1661)
        );

 
    UMUL_1662 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1662),
            data_im_in => first_stage_im_out(1662),
            re_multiplicator => "0000001011000000", --- 0.04296875 + j0.999084472656
            im_multiplicator => "0011111111110001",
            data_re_out => mul_re_out(1662),
            data_im_out => mul_im_out(1662)
        );

 
    UMUL_1663 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1663),
            data_im_in => first_stage_im_out(1663),
            re_multiplicator => "0000011110100100", --- 0.119384765625 + j0.992858886719
            im_multiplicator => "0011111110001011",
            data_re_out => mul_re_out(1663),
            data_im_out => mul_im_out(1663)
        );

 
    UMUL_1664 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1664),
            data_im_in => first_stage_im_out(1664),
            data_re_out => mul_re_out(1664),
            data_im_out => mul_im_out(1664)
        );

 
    UMUL_1665 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1665),
            data_im_in => first_stage_im_out(1665),
            re_multiplicator => "0011111111001100", --- 0.996826171875 + j-0.0797119140625
            im_multiplicator => "1111101011100110",
            data_re_out => mul_re_out(1665),
            data_im_out => mul_im_out(1665)
        );

 
    UMUL_1666 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1666),
            data_im_in => first_stage_im_out(1666),
            re_multiplicator => "0011111100110000", --- 0.9873046875 + j-0.158874511719
            im_multiplicator => "1111010111010101",
            data_re_out => mul_re_out(1666),
            data_im_out => mul_im_out(1666)
        );

 
    UMUL_1667 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1667),
            data_im_in => first_stage_im_out(1667),
            re_multiplicator => "0011111000101101", --- 0.971496582031 + j-0.236999511719
            im_multiplicator => "1111000011010101",
            data_re_out => mul_re_out(1667),
            data_im_out => mul_im_out(1667)
        );

 
    UMUL_1668 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1668),
            data_im_in => first_stage_im_out(1668),
            re_multiplicator => "0011110011000101", --- 0.949523925781 + j-0.313659667969
            im_multiplicator => "1110101111101101",
            data_re_out => mul_re_out(1668),
            data_im_out => mul_im_out(1668)
        );

 
    UMUL_1669 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1669),
            data_im_in => first_stage_im_out(1669),
            re_multiplicator => "0011101011111010", --- 0.921508789062 + j-0.388366699219
            im_multiplicator => "1110011100100101",
            data_re_out => mul_re_out(1669),
            data_im_out => mul_im_out(1669)
        );

 
    UMUL_1670 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1670),
            data_im_in => first_stage_im_out(1670),
            re_multiplicator => "0011100011001111", --- 0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(1670),
            data_im_out => mul_im_out(1670)
        );

 
    UMUL_1671 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1671),
            data_im_in => first_stage_im_out(1671),
            re_multiplicator => "0011011001001000", --- 0.84814453125 + j-0.52978515625
            im_multiplicator => "1101111000011000",
            data_re_out => mul_re_out(1671),
            data_im_out => mul_im_out(1671)
        );

 
    UMUL_1672 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1672),
            data_im_in => first_stage_im_out(1672),
            re_multiplicator => "0011001101101000", --- 0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(1672),
            data_im_out => mul_im_out(1672)
        );

 
    UMUL_1673 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1673),
            data_im_in => first_stage_im_out(1673),
            re_multiplicator => "0011000000110100", --- 0.753173828125 + j-0.657836914062
            im_multiplicator => "1101010111100110",
            data_re_out => mul_re_out(1673),
            data_im_out => mul_im_out(1673)
        );

 
    UMUL_1674 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1674),
            data_im_in => first_stage_im_out(1674),
            re_multiplicator => "0010110010110010", --- 0.698364257812 + j-0.715759277344
            im_multiplicator => "1101001000110001",
            data_re_out => mul_re_out(1674),
            data_im_out => mul_im_out(1674)
        );

 
    UMUL_1675 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1675),
            data_im_in => first_stage_im_out(1675),
            re_multiplicator => "0010100011100111", --- 0.639099121094 + j-0.769104003906
            im_multiplicator => "1100111011000111",
            data_re_out => mul_re_out(1675),
            data_im_out => mul_im_out(1675)
        );

 
    UMUL_1676 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1676),
            data_im_in => first_stage_im_out(1676),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j-0.817565917969
            im_multiplicator => "1100101110101101",
            data_re_out => mul_re_out(1676),
            data_im_out => mul_im_out(1676)
        );

 
    UMUL_1677 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1677),
            data_im_in => first_stage_im_out(1677),
            re_multiplicator => "0010000010010001", --- 0.508850097656 + j-0.86083984375
            im_multiplicator => "1100100011101000",
            data_re_out => mul_re_out(1677),
            data_im_out => mul_im_out(1677)
        );

 
    UMUL_1678 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1678),
            data_im_in => first_stage_im_out(1678),
            re_multiplicator => "0001110000010010", --- 0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(1678),
            data_im_out => mul_im_out(1678)
        );

 
    UMUL_1679 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1679),
            data_im_in => first_stage_im_out(1679),
            re_multiplicator => "0001011101100110", --- 0.365600585938 + j-0.930786132812
            im_multiplicator => "1100010001101110",
            data_re_out => mul_re_out(1679),
            data_im_out => mul_im_out(1679)
        );

 
    UMUL_1680 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1680),
            data_im_in => first_stage_im_out(1680),
            re_multiplicator => "0001001010010100", --- 0.290283203125 + j-0.956970214844
            im_multiplicator => "1100001011000001",
            data_re_out => mul_re_out(1680),
            data_im_out => mul_im_out(1680)
        );

 
    UMUL_1681 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1681),
            data_im_in => first_stage_im_out(1681),
            re_multiplicator => "0000110110100100", --- 0.213134765625 + j-0.97705078125
            im_multiplicator => "1100000101111000",
            data_re_out => mul_re_out(1681),
            data_im_out => mul_im_out(1681)
        );

 
    UMUL_1682 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1682),
            data_im_in => first_stage_im_out(1682),
            re_multiplicator => "0000100010011101", --- 0.134582519531 + j-0.990905761719
            im_multiplicator => "1100000010010101",
            data_re_out => mul_re_out(1682),
            data_im_out => mul_im_out(1682)
        );

 
    UMUL_1683 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1683),
            data_im_in => first_stage_im_out(1683),
            re_multiplicator => "0000001110001000", --- 0.05517578125 + j-0.998474121094
            im_multiplicator => "1100000000011001",
            data_re_out => mul_re_out(1683),
            data_im_out => mul_im_out(1683)
        );

 
    UMUL_1684 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1684),
            data_im_in => first_stage_im_out(1684),
            re_multiplicator => "1111111001101110", --- -0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(1684),
            data_im_out => mul_im_out(1684)
        );

 
    UMUL_1685 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1685),
            data_im_in => first_stage_im_out(1685),
            re_multiplicator => "1111100101010110", --- -0.104125976562 + j-0.994567871094
            im_multiplicator => "1100000001011001",
            data_re_out => mul_re_out(1685),
            data_im_out => mul_im_out(1685)
        );

 
    UMUL_1686 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1686),
            data_im_in => first_stage_im_out(1686),
            re_multiplicator => "1111010001001001", --- -0.183044433594 + j-0.983093261719
            im_multiplicator => "1100000100010101",
            data_re_out => mul_re_out(1686),
            data_im_out => mul_im_out(1686)
        );

 
    UMUL_1687 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1687),
            data_im_in => first_stage_im_out(1687),
            re_multiplicator => "1110111101001111", --- -0.260803222656 + j-0.965393066406
            im_multiplicator => "1100001000110111",
            data_re_out => mul_re_out(1687),
            data_im_out => mul_im_out(1687)
        );

 
    UMUL_1688 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1688),
            data_im_in => first_stage_im_out(1688),
            re_multiplicator => "1110101001110000", --- -0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(1688),
            data_im_out => mul_im_out(1688)
        );

 
    UMUL_1689 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1689),
            data_im_in => first_stage_im_out(1689),
            re_multiplicator => "1110010110110101", --- -0.410827636719 + j-0.911682128906
            im_multiplicator => "1100010110100111",
            data_re_out => mul_re_out(1689),
            data_im_out => mul_im_out(1689)
        );

 
    UMUL_1690 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1690),
            data_im_in => first_stage_im_out(1690),
            re_multiplicator => "1110000100100100", --- -0.482177734375 + j-0.876098632812
            im_multiplicator => "1100011111101110",
            data_re_out => mul_re_out(1690),
            data_im_out => mul_im_out(1690)
        );

 
    UMUL_1691 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1691),
            data_im_in => first_stage_im_out(1691),
            re_multiplicator => "1101110011000101", --- -0.550476074219 + j-0.834838867188
            im_multiplicator => "1100101010010010",
            data_re_out => mul_re_out(1691),
            data_im_out => mul_im_out(1691)
        );

 
    UMUL_1692 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1692),
            data_im_in => first_stage_im_out(1692),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j-0.788330078125
            im_multiplicator => "1100110110001100",
            data_re_out => mul_re_out(1692),
            data_im_out => mul_im_out(1692)
        );

 
    UMUL_1693 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1693),
            data_im_in => first_stage_im_out(1693),
            re_multiplicator => "1101010010111011", --- -0.676086425781 + j-0.73681640625
            im_multiplicator => "1101000011011000",
            data_re_out => mul_re_out(1693),
            data_im_out => mul_im_out(1693)
        );

 
    UMUL_1694 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1694),
            data_im_in => first_stage_im_out(1694),
            re_multiplicator => "1101000100011100", --- -0.732666015625 + j-0.680603027344
            im_multiplicator => "1101010001110001",
            data_re_out => mul_re_out(1694),
            data_im_out => mul_im_out(1694)
        );

 
    UMUL_1695 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1695),
            data_im_in => first_stage_im_out(1695),
            re_multiplicator => "1100110111001010", --- -0.784545898438 + j-0.620056152344
            im_multiplicator => "1101100001010001",
            data_re_out => mul_re_out(1695),
            data_im_out => mul_im_out(1695)
        );

 
    UMUL_1696 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1696),
            data_im_in => first_stage_im_out(1696),
            re_multiplicator => "1100101011001001", --- -0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(1696),
            data_im_out => mul_im_out(1696)
        );

 
    UMUL_1697 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1697),
            data_im_in => first_stage_im_out(1697),
            re_multiplicator => "1100100000011111", --- -0.873107910156 + j-0.487548828125
            im_multiplicator => "1110000011001100",
            data_re_out => mul_re_out(1697),
            data_im_out => mul_im_out(1697)
        );

 
    UMUL_1698 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1698),
            data_im_in => first_stage_im_out(1698),
            re_multiplicator => "1100010111010000", --- -0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(1698),
            data_im_out => mul_im_out(1698)
        );

 
    UMUL_1699 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1699),
            data_im_in => first_stage_im_out(1699),
            re_multiplicator => "1100001111100000", --- -0.939453125 + j-0.342651367188
            im_multiplicator => "1110101000010010",
            data_re_out => mul_re_out(1699),
            data_im_out => mul_im_out(1699)
        );

 
    UMUL_1700 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1700),
            data_im_in => first_stage_im_out(1700),
            re_multiplicator => "1100001001010001", --- -0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(1700),
            data_im_out => mul_im_out(1700)
        );

 
    UMUL_1701 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1701),
            data_im_in => first_stage_im_out(1701),
            re_multiplicator => "1100000100101000", --- -0.98193359375 + j-0.189086914062
            im_multiplicator => "1111001111100110",
            data_re_out => mul_re_out(1701),
            data_im_out => mul_im_out(1701)
        );

 
    UMUL_1702 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1702),
            data_im_in => first_stage_im_out(1702),
            re_multiplicator => "1100000001100100", --- -0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(1702),
            data_im_out => mul_im_out(1702)
        );

 
    UMUL_1703 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1703),
            data_im_in => first_stage_im_out(1703),
            re_multiplicator => "1100000000001000", --- -0.99951171875 + j-0.0307006835938
            im_multiplicator => "1111111000001001",
            data_re_out => mul_re_out(1703),
            data_im_out => mul_im_out(1703)
        );

 
    UMUL_1704 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1704),
            data_im_in => first_stage_im_out(1704),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j0.049072265625
            im_multiplicator => "0000001100100100",
            data_re_out => mul_re_out(1704),
            data_im_out => mul_im_out(1704)
        );

 
    UMUL_1705 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1705),
            data_im_in => first_stage_im_out(1705),
            re_multiplicator => "1100000010001000", --- -0.99169921875 + j0.128479003906
            im_multiplicator => "0000100000111001",
            data_re_out => mul_re_out(1705),
            data_im_out => mul_im_out(1705)
        );

 
    UMUL_1706 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1706),
            data_im_in => first_stage_im_out(1706),
            re_multiplicator => "1100000101100011", --- -0.978332519531 + j0.207092285156
            im_multiplicator => "0000110101000001",
            data_re_out => mul_re_out(1706),
            data_im_out => mul_im_out(1706)
        );

 
    UMUL_1707 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1707),
            data_im_in => first_stage_im_out(1707),
            re_multiplicator => "1100001010100101", --- -0.958679199219 + j0.284423828125
            im_multiplicator => "0001001000110100",
            data_re_out => mul_re_out(1707),
            data_im_out => mul_im_out(1707)
        );

 
    UMUL_1708 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1708),
            data_im_in => first_stage_im_out(1708),
            re_multiplicator => "1100010001001010", --- -0.932983398438 + j0.359924316406
            im_multiplicator => "0001011100001001",
            data_re_out => mul_re_out(1708),
            data_im_out => mul_im_out(1708)
        );

 
    UMUL_1709 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1709),
            data_im_in => first_stage_im_out(1709),
            re_multiplicator => "1100011001010000", --- -0.9013671875 + j0.43310546875
            im_multiplicator => "0001101110111000",
            data_re_out => mul_re_out(1709),
            data_im_out => mul_im_out(1709)
        );

 
    UMUL_1710 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1710),
            data_im_in => first_stage_im_out(1710),
            re_multiplicator => "1100100010110101", --- -0.863952636719 + j0.503540039062
            im_multiplicator => "0010000000111010",
            data_re_out => mul_re_out(1710),
            data_im_out => mul_im_out(1710)
        );

 
    UMUL_1711 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1711),
            data_im_in => first_stage_im_out(1711),
            re_multiplicator => "1100101101110011", --- -0.821105957031 + j0.57080078125
            im_multiplicator => "0010010010001000",
            data_re_out => mul_re_out(1711),
            data_im_out => mul_im_out(1711)
        );

 
    UMUL_1712 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1712),
            data_im_in => first_stage_im_out(1712),
            re_multiplicator => "1100111010000111", --- -0.773010253906 + j0.634399414062
            im_multiplicator => "0010100010011010",
            data_re_out => mul_re_out(1712),
            data_im_out => mul_im_out(1712)
        );

 
    UMUL_1713 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1713),
            data_im_in => first_stage_im_out(1713),
            re_multiplicator => "1101000111101011", --- -0.720031738281 + j0.693969726562
            im_multiplicator => "0010110001101010",
            data_re_out => mul_re_out(1713),
            data_im_out => mul_im_out(1713)
        );

 
    UMUL_1714 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1714),
            data_im_in => first_stage_im_out(1714),
            re_multiplicator => "1101010110011011", --- -0.662414550781 + j0.749145507812
            im_multiplicator => "0010111111110010",
            data_re_out => mul_re_out(1714),
            data_im_out => mul_im_out(1714)
        );

 
    UMUL_1715 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1715),
            data_im_in => first_stage_im_out(1715),
            re_multiplicator => "1101100110001111", --- -0.600646972656 + j0.799560546875
            im_multiplicator => "0011001100101100",
            data_re_out => mul_re_out(1715),
            data_im_out => mul_im_out(1715)
        );

 
    UMUL_1716 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1716),
            data_im_in => first_stage_im_out(1716),
            re_multiplicator => "1101110111000011", --- -0.534973144531 + j0.844848632812
            im_multiplicator => "0011011000010010",
            data_re_out => mul_re_out(1716),
            data_im_out => mul_im_out(1716)
        );

 
    UMUL_1717 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1717),
            data_im_in => first_stage_im_out(1717),
            re_multiplicator => "1110001000101101", --- -0.466003417969 + j0.884826660156
            im_multiplicator => "0011100010100001",
            data_re_out => mul_re_out(1717),
            data_im_out => mul_im_out(1717)
        );

 
    UMUL_1718 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1718),
            data_im_in => first_stage_im_out(1718),
            re_multiplicator => "1110011011001001", --- -0.393981933594 + j0.919128417969
            im_multiplicator => "0011101011010011",
            data_re_out => mul_re_out(1718),
            data_im_out => mul_im_out(1718)
        );

 
    UMUL_1719 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1719),
            data_im_in => first_stage_im_out(1719),
            re_multiplicator => "1110101110001101", --- -0.319519042969 + j0.947570800781
            im_multiplicator => "0011110010100101",
            data_re_out => mul_re_out(1719),
            data_im_out => mul_im_out(1719)
        );

 
    UMUL_1720 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1720),
            data_im_in => first_stage_im_out(1720),
            re_multiplicator => "1111000001110011", --- -0.242980957031 + j0.970031738281
            im_multiplicator => "0011111000010101",
            data_re_out => mul_re_out(1720),
            data_im_out => mul_im_out(1720)
        );

 
    UMUL_1721 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1721),
            data_im_in => first_stage_im_out(1721),
            re_multiplicator => "1111010101110010", --- -0.164916992188 + j0.986328125
            im_multiplicator => "0011111100100000",
            data_re_out => mul_re_out(1721),
            data_im_out => mul_im_out(1721)
        );

 
    UMUL_1722 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1722),
            data_im_in => first_stage_im_out(1722),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j0.996337890625
            im_multiplicator => "0011111111000100",
            data_re_out => mul_re_out(1722),
            data_im_out => mul_im_out(1722)
        );

 
    UMUL_1723 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1723),
            data_im_in => first_stage_im_out(1723),
            re_multiplicator => "1111111110011011", --- -0.00616455078125 + j1.0
            im_multiplicator => "0100000000000000",
            data_re_out => mul_re_out(1723),
            data_im_out => mul_im_out(1723)
        );

 
    UMUL_1724 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1724),
            data_im_in => first_stage_im_out(1724),
            re_multiplicator => "0000010010110101", --- 0.0735473632812 + j0.997314453125
            im_multiplicator => "0011111111010100",
            data_re_out => mul_re_out(1724),
            data_im_out => mul_im_out(1724)
        );

 
    UMUL_1725 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1725),
            data_im_in => first_stage_im_out(1725),
            re_multiplicator => "0000100111000111", --- 0.152770996094 + j0.98828125
            im_multiplicator => "0011111101000000",
            data_re_out => mul_re_out(1725),
            data_im_out => mul_im_out(1725)
        );

 
    UMUL_1726 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1726),
            data_im_in => first_stage_im_out(1726),
            re_multiplicator => "0000111011001010", --- 0.231079101562 + j0.972961425781
            im_multiplicator => "0011111001000101",
            data_re_out => mul_re_out(1726),
            data_im_out => mul_im_out(1726)
        );

 
    UMUL_1727 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1727),
            data_im_in => first_stage_im_out(1727),
            re_multiplicator => "0001001110110100", --- 0.307861328125 + j0.951416015625
            im_multiplicator => "0011110011100100",
            data_re_out => mul_re_out(1727),
            data_im_out => mul_im_out(1727)
        );

 
    UMUL_1728 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1728),
            data_im_in => first_stage_im_out(1728),
            data_re_out => mul_re_out(1728),
            data_im_out => mul_im_out(1728)
        );

 
    UMUL_1729 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1729),
            data_im_in => first_stage_im_out(1729),
            re_multiplicator => "0011111111001000", --- 0.99658203125 + j-0.082763671875
            im_multiplicator => "1111101010110100",
            data_re_out => mul_re_out(1729),
            data_im_out => mul_im_out(1729)
        );

 
    UMUL_1730 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1730),
            data_im_in => first_stage_im_out(1730),
            re_multiplicator => "0011111100100000", --- 0.986328125 + j-0.164916992188
            im_multiplicator => "1111010101110010",
            data_re_out => mul_re_out(1730),
            data_im_out => mul_im_out(1730)
        );

 
    UMUL_1731 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1731),
            data_im_in => first_stage_im_out(1731),
            re_multiplicator => "0011111000001001", --- 0.969299316406 + j-0.245971679688
            im_multiplicator => "1111000001000010",
            data_re_out => mul_re_out(1731),
            data_im_out => mul_im_out(1731)
        );

 
    UMUL_1732 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1732),
            data_im_in => first_stage_im_out(1732),
            re_multiplicator => "0011110010000101", --- 0.945617675781 + j-0.325317382812
            im_multiplicator => "1110101100101110",
            data_re_out => mul_re_out(1732),
            data_im_out => mul_im_out(1732)
        );

 
    UMUL_1733 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1733),
            data_im_in => first_stage_im_out(1733),
            re_multiplicator => "0011101010010111", --- 0.915466308594 + j-0.402404785156
            im_multiplicator => "1110011000111111",
            data_re_out => mul_re_out(1733),
            data_im_out => mul_im_out(1733)
        );

 
    UMUL_1734 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1734),
            data_im_in => first_stage_im_out(1734),
            re_multiplicator => "0011100001000010", --- 0.879028320312 + j-0.476806640625
            im_multiplicator => "1110000101111100",
            data_re_out => mul_re_out(1734),
            data_im_out => mul_im_out(1734)
        );

 
    UMUL_1735 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1735),
            data_im_in => first_stage_im_out(1735),
            re_multiplicator => "0011010110001010", --- 0.836547851562 + j-0.547912597656
            im_multiplicator => "1101110011101111",
            data_re_out => mul_re_out(1735),
            data_im_out => mul_im_out(1735)
        );

 
    UMUL_1736 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1736),
            data_im_in => first_stage_im_out(1736),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(1736),
            data_im_out => mul_im_out(1736)
        );

 
    UMUL_1737 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1737),
            data_im_in => first_stage_im_out(1737),
            re_multiplicator => "0010111100000110", --- 0.734741210938 + j-0.678344726562
            im_multiplicator => "1101010010010110",
            data_re_out => mul_re_out(1737),
            data_im_out => mul_im_out(1737)
        );

 
    UMUL_1738 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1738),
            data_im_in => first_stage_im_out(1738),
            re_multiplicator => "0010101101000101", --- 0.676086425781 + j-0.73681640625
            im_multiplicator => "1101000011011000",
            data_re_out => mul_re_out(1738),
            data_im_out => mul_im_out(1738)
        );

 
    UMUL_1739 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1739),
            data_im_in => first_stage_im_out(1739),
            re_multiplicator => "0010011100111000", --- 0.61279296875 + j-0.790222167969
            im_multiplicator => "1100110101101101",
            data_re_out => mul_re_out(1739),
            data_im_out => mul_im_out(1739)
        );

 
    UMUL_1740 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1740),
            data_im_in => first_stage_im_out(1740),
            re_multiplicator => "0010001011100111", --- 0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(1740),
            data_im_out => mul_im_out(1740)
        );

 
    UMUL_1741 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1741),
            data_im_in => first_stage_im_out(1741),
            re_multiplicator => "0001111001011000", --- 0.47412109375 + j-0.880493164062
            im_multiplicator => "1100011110100110",
            data_re_out => mul_re_out(1741),
            data_im_out => mul_im_out(1741)
        );

 
    UMUL_1742 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1742),
            data_im_in => first_stage_im_out(1742),
            re_multiplicator => "0001100110010011", --- 0.399597167969 + j-0.916687011719
            im_multiplicator => "1100010101010101",
            data_re_out => mul_re_out(1742),
            data_im_out => mul_im_out(1742)
        );

 
    UMUL_1743 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1743),
            data_im_in => first_stage_im_out(1743),
            re_multiplicator => "0001010010100010", --- 0.322387695312 + j-0.946594238281
            im_multiplicator => "1100001101101011",
            data_re_out => mul_re_out(1743),
            data_im_out => mul_im_out(1743)
        );

 
    UMUL_1744 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1744),
            data_im_in => first_stage_im_out(1744),
            re_multiplicator => "0000111110001101", --- 0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(1744),
            data_im_out => mul_im_out(1744)
        );

 
    UMUL_1745 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1745),
            data_im_in => first_stage_im_out(1745),
            re_multiplicator => "0000101001011100", --- 0.161865234375 + j-0.98681640625
            im_multiplicator => "1100000011011000",
            data_re_out => mul_re_out(1745),
            data_im_out => mul_im_out(1745)
        );

 
    UMUL_1746 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1746),
            data_im_in => first_stage_im_out(1746),
            re_multiplicator => "0000010100011010", --- 0.0797119140625 + j-0.996826171875
            im_multiplicator => "1100000000110100",
            data_re_out => mul_re_out(1746),
            data_im_out => mul_im_out(1746)
        );

 
    UMUL_1747 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1747),
            data_im_in => first_stage_im_out(1747),
            re_multiplicator => "1111111111001110", --- -0.0030517578125 + j-1.0
            im_multiplicator => "1100000000000000",
            data_re_out => mul_re_out(1747),
            data_im_out => mul_im_out(1747)
        );

 
    UMUL_1748 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1748),
            data_im_in => first_stage_im_out(1748),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(1748),
            data_im_out => mul_im_out(1748)
        );

 
    UMUL_1749 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1749),
            data_im_in => first_stage_im_out(1749),
            re_multiplicator => "1111010101000000", --- -0.16796875 + j-0.985778808594
            im_multiplicator => "1100000011101001",
            data_re_out => mul_re_out(1749),
            data_im_out => mul_im_out(1749)
        );

 
    UMUL_1750 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1750),
            data_im_in => first_stage_im_out(1750),
            re_multiplicator => "1111000000010010", --- -0.248901367188 + j-0.968505859375
            im_multiplicator => "1100001000000100",
            data_re_out => mul_re_out(1750),
            data_im_out => mul_im_out(1750)
        );

 
    UMUL_1751 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1751),
            data_im_in => first_stage_im_out(1751),
            re_multiplicator => "1110101011111111", --- -0.328186035156 + j-0.944580078125
            im_multiplicator => "1100001110001100",
            data_re_out => mul_re_out(1751),
            data_im_out => mul_im_out(1751)
        );

 
    UMUL_1752 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1752),
            data_im_in => first_stage_im_out(1752),
            re_multiplicator => "1110011000010001", --- -0.405212402344 + j-0.914184570312
            im_multiplicator => "1100010101111110",
            data_re_out => mul_re_out(1752),
            data_im_out => mul_im_out(1752)
        );

 
    UMUL_1753 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1753),
            data_im_in => first_stage_im_out(1753),
            re_multiplicator => "1110000101010000", --- -0.4794921875 + j-0.877563476562
            im_multiplicator => "1100011111010110",
            data_re_out => mul_re_out(1753),
            data_im_out => mul_im_out(1753)
        );

 
    UMUL_1754 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1754),
            data_im_in => first_stage_im_out(1754),
            re_multiplicator => "1101110011000101", --- -0.550476074219 + j-0.834838867188
            im_multiplicator => "1100101010010010",
            data_re_out => mul_re_out(1754),
            data_im_out => mul_im_out(1754)
        );

 
    UMUL_1755 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1755),
            data_im_in => first_stage_im_out(1755),
            re_multiplicator => "1101100001111000", --- -0.61767578125 + j-0.786437988281
            im_multiplicator => "1100110110101011",
            data_re_out => mul_re_out(1755),
            data_im_out => mul_im_out(1755)
        );

 
    UMUL_1756 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1756),
            data_im_in => first_stage_im_out(1756),
            re_multiplicator => "1101010001110001", --- -0.680603027344 + j-0.732666015625
            im_multiplicator => "1101000100011100",
            data_re_out => mul_re_out(1756),
            data_im_out => mul_im_out(1756)
        );

 
    UMUL_1757 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1757),
            data_im_in => first_stage_im_out(1757),
            re_multiplicator => "1101000010110110", --- -0.738891601562 + j-0.673828125
            im_multiplicator => "1101010011100000",
            data_re_out => mul_re_out(1757),
            data_im_out => mul_im_out(1757)
        );

 
    UMUL_1758 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1758),
            data_im_in => first_stage_im_out(1758),
            re_multiplicator => "1100110101001110", --- -0.792114257812 + j-0.610412597656
            im_multiplicator => "1101100011101111",
            data_re_out => mul_re_out(1758),
            data_im_out => mul_im_out(1758)
        );

 
    UMUL_1759 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1759),
            data_im_in => first_stage_im_out(1759),
            re_multiplicator => "1100101000111111", --- -0.839904785156 + j-0.542724609375
            im_multiplicator => "1101110101000100",
            data_re_out => mul_re_out(1759),
            data_im_out => mul_im_out(1759)
        );

 
    UMUL_1760 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1760),
            data_im_in => first_stage_im_out(1760),
            re_multiplicator => "1100011110001111", --- -0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(1760),
            data_im_out => mul_im_out(1760)
        );

 
    UMUL_1761 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1761),
            data_im_in => first_stage_im_out(1761),
            re_multiplicator => "1100010101000001", --- -0.917907714844 + j-0.396789550781
            im_multiplicator => "1110011010011011",
            data_re_out => mul_re_out(1761),
            data_im_out => mul_im_out(1761)
        );

 
    UMUL_1762 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1762),
            data_im_in => first_stage_im_out(1762),
            re_multiplicator => "1100001101011011", --- -0.947570800781 + j-0.319519042969
            im_multiplicator => "1110101110001101",
            data_re_out => mul_re_out(1762),
            data_im_out => mul_im_out(1762)
        );

 
    UMUL_1763 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1763),
            data_im_in => first_stage_im_out(1763),
            re_multiplicator => "1100000111011111", --- -0.970764160156 + j-0.239990234375
            im_multiplicator => "1111000010100100",
            data_re_out => mul_re_out(1763),
            data_im_out => mul_im_out(1763)
        );

 
    UMUL_1764 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1764),
            data_im_in => first_stage_im_out(1764),
            re_multiplicator => "1100000011010000", --- -0.9873046875 + j-0.158874511719
            im_multiplicator => "1111010111010101",
            data_re_out => mul_re_out(1764),
            data_im_out => mul_im_out(1764)
        );

 
    UMUL_1765 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1765),
            data_im_in => first_stage_im_out(1765),
            re_multiplicator => "1100000000110000", --- -0.9970703125 + j-0.0765991210938
            im_multiplicator => "1111101100011001",
            data_re_out => mul_re_out(1765),
            data_im_out => mul_im_out(1765)
        );

 
    UMUL_1766 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1766),
            data_im_in => first_stage_im_out(1766),
            re_multiplicator => "1100000000000000", --- -1.0 + j0.00616455078125
            im_multiplicator => "0000000001100101",
            data_re_out => mul_re_out(1766),
            data_im_out => mul_im_out(1766)
        );

 
    UMUL_1767 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1767),
            data_im_in => first_stage_im_out(1767),
            re_multiplicator => "1100000001000001", --- -0.996032714844 + j0.0888671875
            im_multiplicator => "0000010110110000",
            data_re_out => mul_re_out(1767),
            data_im_out => mul_im_out(1767)
        );

 
    UMUL_1768 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1768),
            data_im_in => first_stage_im_out(1768),
            re_multiplicator => "1100000011110001", --- -0.985290527344 + j0.170959472656
            im_multiplicator => "0000101011110001",
            data_re_out => mul_re_out(1768),
            data_im_out => mul_im_out(1768)
        );

 
    UMUL_1769 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1769),
            data_im_in => first_stage_im_out(1769),
            re_multiplicator => "1100001000010000", --- -0.9677734375 + j0.251892089844
            im_multiplicator => "0001000000011111",
            data_re_out => mul_re_out(1769),
            data_im_out => mul_im_out(1769)
        );

 
    UMUL_1770 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1770),
            data_im_in => first_stage_im_out(1770),
            re_multiplicator => "1100001110011100", --- -0.943603515625 + j0.331115722656
            im_multiplicator => "0001010100110001",
            data_re_out => mul_re_out(1770),
            data_im_out => mul_im_out(1770)
        );

 
    UMUL_1771 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1771),
            data_im_in => first_stage_im_out(1771),
            re_multiplicator => "1100010110010010", --- -0.912963867188 + j0.408020019531
            im_multiplicator => "0001101000011101",
            data_re_out => mul_re_out(1771),
            data_im_out => mul_im_out(1771)
        );

 
    UMUL_1772 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1772),
            data_im_in => first_stage_im_out(1772),
            re_multiplicator => "1100011111101110", --- -0.876098632812 + j0.482177734375
            im_multiplicator => "0001111011011100",
            data_re_out => mul_re_out(1772),
            data_im_out => mul_im_out(1772)
        );

 
    UMUL_1773 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1773),
            data_im_in => first_stage_im_out(1773),
            re_multiplicator => "1100101010101101", --- -0.833190917969 + j0.553039550781
            im_multiplicator => "0010001101100101",
            data_re_out => mul_re_out(1773),
            data_im_out => mul_im_out(1773)
        );

 
    UMUL_1774 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1774),
            data_im_in => first_stage_im_out(1774),
            re_multiplicator => "1100110111001010", --- -0.784545898438 + j0.620056152344
            im_multiplicator => "0010011110101111",
            data_re_out => mul_re_out(1774),
            data_im_out => mul_im_out(1774)
        );

 
    UMUL_1775 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1775),
            data_im_in => first_stage_im_out(1775),
            re_multiplicator => "1101000100111110", --- -0.730590820312 + j0.682861328125
            im_multiplicator => "0010101110110100",
            data_re_out => mul_re_out(1775),
            data_im_out => mul_im_out(1775)
        );

 
    UMUL_1776 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1776),
            data_im_in => first_stage_im_out(1776),
            re_multiplicator => "1101010100000101", --- -0.671569824219 + j0.740966796875
            im_multiplicator => "0010111101101100",
            data_re_out => mul_re_out(1776),
            data_im_out => mul_im_out(1776)
        );

 
    UMUL_1777 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1777),
            data_im_in => first_stage_im_out(1777),
            re_multiplicator => "1101100100010111", --- -0.607971191406 + j0.7939453125
            im_multiplicator => "0011001011010000",
            data_re_out => mul_re_out(1777),
            data_im_out => mul_im_out(1777)
        );

 
    UMUL_1778 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1778),
            data_im_in => first_stage_im_out(1778),
            re_multiplicator => "1101110101101110", --- -0.540161132812 + j0.841552734375
            im_multiplicator => "0011010111011100",
            data_re_out => mul_re_out(1778),
            data_im_out => mul_im_out(1778)
        );

 
    UMUL_1779 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1779),
            data_im_in => first_stage_im_out(1779),
            re_multiplicator => "1110001000000001", --- -0.468688964844 + j0.883361816406
            im_multiplicator => "0011100010001001",
            data_re_out => mul_re_out(1779),
            data_im_out => mul_im_out(1779)
        );

 
    UMUL_1780 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1780),
            data_im_in => first_stage_im_out(1780),
            re_multiplicator => "1110011011001001", --- -0.393981933594 + j0.919128417969
            im_multiplicator => "0011101011010011",
            data_re_out => mul_re_out(1780),
            data_im_out => mul_im_out(1780)
        );

 
    UMUL_1781 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1781),
            data_im_in => first_stage_im_out(1781),
            re_multiplicator => "1110101110111101", --- -0.316589355469 + j0.948547363281
            im_multiplicator => "0011110010110101",
            data_re_out => mul_re_out(1781),
            data_im_out => mul_im_out(1781)
        );

 
    UMUL_1782 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1782),
            data_im_in => first_stage_im_out(1782),
            re_multiplicator => "1111000011010101", --- -0.236999511719 + j0.971496582031
            im_multiplicator => "0011111000101101",
            data_re_out => mul_re_out(1782),
            data_im_out => mul_im_out(1782)
        );

 
    UMUL_1783 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1783),
            data_im_in => first_stage_im_out(1783),
            re_multiplicator => "1111011000000111", --- -0.155822753906 + j0.98779296875
            im_multiplicator => "0011111100111000",
            data_re_out => mul_re_out(1783),
            data_im_out => mul_im_out(1783)
        );

 
    UMUL_1784 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1784),
            data_im_in => first_stage_im_out(1784),
            re_multiplicator => "1111101101001011", --- -0.0735473632812 + j0.997314453125
            im_multiplicator => "0011111111010100",
            data_re_out => mul_re_out(1784),
            data_im_out => mul_im_out(1784)
        );

 
    UMUL_1785 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1785),
            data_im_in => first_stage_im_out(1785),
            re_multiplicator => "0000000010010111", --- 0.00921630859375 + j0.999938964844
            im_multiplicator => "0011111111111111",
            data_re_out => mul_re_out(1785),
            data_im_out => mul_im_out(1785)
        );

 
    UMUL_1786 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1786),
            data_im_in => first_stage_im_out(1786),
            re_multiplicator => "0000010111100010", --- 0.0919189453125 + j0.995788574219
            im_multiplicator => "0011111110111011",
            data_re_out => mul_re_out(1786),
            data_im_out => mul_im_out(1786)
        );

 
    UMUL_1787 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1787),
            data_im_in => first_stage_im_out(1787),
            re_multiplicator => "0000101100100011", --- 0.174011230469 + j0.984741210938
            im_multiplicator => "0011111100000110",
            data_re_out => mul_re_out(1787),
            data_im_out => mul_im_out(1787)
        );

 
    UMUL_1788 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1788),
            data_im_in => first_stage_im_out(1788),
            re_multiplicator => "0001000001010000", --- 0.2548828125 + j0.966979980469
            im_multiplicator => "0011110111100011",
            data_re_out => mul_re_out(1788),
            data_im_out => mul_im_out(1788)
        );

 
    UMUL_1789 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1789),
            data_im_in => first_stage_im_out(1789),
            re_multiplicator => "0001010101100000", --- 0.333984375 + j0.942565917969
            im_multiplicator => "0011110001010011",
            data_re_out => mul_re_out(1789),
            data_im_out => mul_im_out(1789)
        );

 
    UMUL_1790 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1790),
            data_im_in => first_stage_im_out(1790),
            re_multiplicator => "0001101001001011", --- 0.410827636719 + j0.911682128906
            im_multiplicator => "0011101001011001",
            data_re_out => mul_re_out(1790),
            data_im_out => mul_im_out(1790)
        );

 
    UMUL_1791 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1791),
            data_im_in => first_stage_im_out(1791),
            re_multiplicator => "0001111100001000", --- 0.48486328125 + j0.874572753906
            im_multiplicator => "0011011111111001",
            data_re_out => mul_re_out(1791),
            data_im_out => mul_im_out(1791)
        );

 
    UMUL_1792 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1792),
            data_im_in => first_stage_im_out(1792),
            data_re_out => mul_re_out(1792),
            data_im_out => mul_im_out(1792)
        );

 
    UMUL_1793 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1793),
            data_im_in => first_stage_im_out(1793),
            re_multiplicator => "0011111111000100", --- 0.996337890625 + j-0.0858154296875
            im_multiplicator => "1111101010000010",
            data_re_out => mul_re_out(1793),
            data_im_out => mul_im_out(1793)
        );

 
    UMUL_1794 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1794),
            data_im_in => first_stage_im_out(1794),
            re_multiplicator => "0011111100001111", --- 0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(1794),
            data_im_out => mul_im_out(1794)
        );

 
    UMUL_1795 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1795),
            data_im_in => first_stage_im_out(1795),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(1795),
            data_im_out => mul_im_out(1795)
        );

 
    UMUL_1796 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1796),
            data_im_in => first_stage_im_out(1796),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(1796),
            data_im_out => mul_im_out(1796)
        );

 
    UMUL_1797 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1797),
            data_im_in => first_stage_im_out(1797),
            re_multiplicator => "0011101000110000", --- 0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(1797),
            data_im_out => mul_im_out(1797)
        );

 
    UMUL_1798 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1798),
            data_im_in => first_stage_im_out(1798),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(1798),
            data_im_out => mul_im_out(1798)
        );

 
    UMUL_1799 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1799),
            data_im_in => first_stage_im_out(1799),
            re_multiplicator => "0011010011000110", --- 0.824584960938 + j-0.565734863281
            im_multiplicator => "1101101111001011",
            data_re_out => mul_re_out(1799),
            data_im_out => mul_im_out(1799)
        );

 
    UMUL_1800 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1800),
            data_im_in => first_stage_im_out(1800),
            re_multiplicator => "0011000101111001", --- 0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(1800),
            data_im_out => mul_im_out(1800)
        );

 
    UMUL_1801 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1801),
            data_im_in => first_stage_im_out(1801),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(1801),
            data_im_out => mul_im_out(1801)
        );

 
    UMUL_1802 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1802),
            data_im_in => first_stage_im_out(1802),
            re_multiplicator => "0010100111001110", --- 0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(1802),
            data_im_out => mul_im_out(1802)
        );

 
    UMUL_1803 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1803),
            data_im_in => first_stage_im_out(1803),
            re_multiplicator => "0010010101111110", --- 0.585815429688 + j-0.810485839844
            im_multiplicator => "1100110000100001",
            data_re_out => mul_re_out(1803),
            data_im_out => mul_im_out(1803)
        );

 
    UMUL_1804 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1804),
            data_im_in => first_stage_im_out(1804),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(1804),
            data_im_out => mul_im_out(1804)
        );

 
    UMUL_1805 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1805),
            data_im_in => first_stage_im_out(1805),
            re_multiplicator => "0001110000010010", --- 0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(1805),
            data_im_out => mul_im_out(1805)
        );

 
    UMUL_1806 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1806),
            data_im_in => first_stage_im_out(1806),
            re_multiplicator => "0001011100001001", --- 0.359924316406 + j-0.932983398438
            im_multiplicator => "1100010001001010",
            data_re_out => mul_re_out(1806),
            data_im_out => mul_im_out(1806)
        );

 
    UMUL_1807 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1807),
            data_im_in => first_stage_im_out(1807),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(1807),
            data_im_out => mul_im_out(1807)
        );

 
    UMUL_1808 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1808),
            data_im_in => first_stage_im_out(1808),
            re_multiplicator => "0000110001111100", --- 0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(1808),
            data_im_out => mul_im_out(1808)
        );

 
    UMUL_1809 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1809),
            data_im_in => first_stage_im_out(1809),
            re_multiplicator => "0000011100001110", --- 0.110229492188 + j-0.993896484375
            im_multiplicator => "1100000001100100",
            data_re_out => mul_re_out(1809),
            data_im_out => mul_im_out(1809)
        );

 
    UMUL_1810 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1810),
            data_im_in => first_stage_im_out(1810),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(1810),
            data_im_out => mul_im_out(1810)
        );

 
    UMUL_1811 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1811),
            data_im_in => first_stage_im_out(1811),
            re_multiplicator => "1111110000010011", --- -0.0613403320312 + j-0.998107910156
            im_multiplicator => "1100000000011111",
            data_re_out => mul_re_out(1811),
            data_im_out => mul_im_out(1811)
        );

 
    UMUL_1812 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1812),
            data_im_in => first_stage_im_out(1812),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(1812),
            data_im_out => mul_im_out(1812)
        );

 
    UMUL_1813 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1813),
            data_im_in => first_stage_im_out(1813),
            re_multiplicator => "1111000100110110", --- -0.231079101562 + j-0.972961425781
            im_multiplicator => "1100000110111011",
            data_re_out => mul_re_out(1813),
            data_im_out => mul_im_out(1813)
        );

 
    UMUL_1814 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1814),
            data_im_in => first_stage_im_out(1814),
            re_multiplicator => "1110101111101101", --- -0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(1814),
            data_im_out => mul_im_out(1814)
        );

 
    UMUL_1815 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1815),
            data_im_in => first_stage_im_out(1815),
            re_multiplicator => "1110011011001001", --- -0.393981933594 + j-0.919128417969
            im_multiplicator => "1100010100101101",
            data_re_out => mul_re_out(1815),
            data_im_out => mul_im_out(1815)
        );

 
    UMUL_1816 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1816),
            data_im_in => first_stage_im_out(1816),
            re_multiplicator => "1110000111010101", --- -0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(1816),
            data_im_out => mul_im_out(1816)
        );

 
    UMUL_1817 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1817),
            data_im_in => first_stage_im_out(1817),
            re_multiplicator => "1101110100011001", --- -0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(1817),
            data_im_out => mul_im_out(1817)
        );

 
    UMUL_1818 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1818),
            data_im_in => first_stage_im_out(1818),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j-0.788330078125
            im_multiplicator => "1100110110001100",
            data_re_out => mul_re_out(1818),
            data_im_out => mul_im_out(1818)
        );

 
    UMUL_1819 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1819),
            data_im_in => first_stage_im_out(1819),
            re_multiplicator => "1101010001110001", --- -0.680603027344 + j-0.732666015625
            im_multiplicator => "1101000100011100",
            data_re_out => mul_re_out(1819),
            data_im_out => mul_im_out(1819)
        );

 
    UMUL_1820 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1820),
            data_im_in => first_stage_im_out(1820),
            re_multiplicator => "1101000010010100", --- -0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(1820),
            data_im_out => mul_im_out(1820)
        );

 
    UMUL_1821 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1821),
            data_im_in => first_stage_im_out(1821),
            re_multiplicator => "1100110100010001", --- -0.795837402344 + j-0.605529785156
            im_multiplicator => "1101100100111111",
            data_re_out => mul_re_out(1821),
            data_im_out => mul_im_out(1821)
        );

 
    UMUL_1822 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1822),
            data_im_in => first_stage_im_out(1822),
            re_multiplicator => "1100100111101110", --- -0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(1822),
            data_im_out => mul_im_out(1822)
        );

 
    UMUL_1823 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1823),
            data_im_in => first_stage_im_out(1823),
            re_multiplicator => "1100011100110001", --- -0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(1823),
            data_im_out => mul_im_out(1823)
        );

 
    UMUL_1824 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1824),
            data_im_in => first_stage_im_out(1824),
            re_multiplicator => "1100010011011111", --- -0.923889160156 + j-0.382690429688
            im_multiplicator => "1110011110000010",
            data_re_out => mul_re_out(1824),
            data_im_out => mul_im_out(1824)
        );

 
    UMUL_1825 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1825),
            data_im_in => first_stage_im_out(1825),
            re_multiplicator => "1100001011111101", --- -0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(1825),
            data_im_out => mul_im_out(1825)
        );

 
    UMUL_1826 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1826),
            data_im_in => first_stage_im_out(1826),
            re_multiplicator => "1100000110001110", --- -0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(1826),
            data_im_out => mul_im_out(1826)
        );

 
    UMUL_1827 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1827),
            data_im_in => first_stage_im_out(1827),
            re_multiplicator => "1100000010010101", --- -0.990905761719 + j-0.134582519531
            im_multiplicator => "1111011101100011",
            data_re_out => mul_re_out(1827),
            data_im_out => mul_im_out(1827)
        );

 
    UMUL_1828 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1828),
            data_im_in => first_stage_im_out(1828),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(1828),
            data_im_out => mul_im_out(1828)
        );

 
    UMUL_1829 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1829),
            data_im_in => first_stage_im_out(1829),
            re_multiplicator => "1100000000001011", --- -0.999328613281 + j0.0368041992188
            im_multiplicator => "0000001001011011",
            data_re_out => mul_re_out(1829),
            data_im_out => mul_im_out(1829)
        );

 
    UMUL_1830 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1830),
            data_im_in => first_stage_im_out(1830),
            re_multiplicator => "1100000001111011", --- -0.992492675781 + j0.122436523438
            im_multiplicator => "0000011111010110",
            data_re_out => mul_re_out(1830),
            data_im_out => mul_im_out(1830)
        );

 
    UMUL_1831 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1831),
            data_im_in => first_stage_im_out(1831),
            re_multiplicator => "1100000101100011", --- -0.978332519531 + j0.207092285156
            im_multiplicator => "0000110101000001",
            data_re_out => mul_re_out(1831),
            data_im_out => mul_im_out(1831)
        );

 
    UMUL_1832 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1832),
            data_im_in => first_stage_im_out(1832),
            re_multiplicator => "1100001011000001", --- -0.956970214844 + j0.290283203125
            im_multiplicator => "0001001010010100",
            data_re_out => mul_re_out(1832),
            data_im_out => mul_im_out(1832)
        );

 
    UMUL_1833 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1833),
            data_im_in => first_stage_im_out(1833),
            re_multiplicator => "1100010010010011", --- -0.928527832031 + j0.371337890625
            im_multiplicator => "0001011111000100",
            data_re_out => mul_re_out(1833),
            data_im_out => mul_im_out(1833)
        );

 
    UMUL_1834 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1834),
            data_im_in => first_stage_im_out(1834),
            re_multiplicator => "1100011011010101", --- -0.893249511719 + j0.449584960938
            im_multiplicator => "0001110011000110",
            data_re_out => mul_re_out(1834),
            data_im_out => mul_im_out(1834)
        );

 
    UMUL_1835 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1835),
            data_im_in => first_stage_im_out(1835),
            re_multiplicator => "1100100110000011", --- -0.851379394531 + j0.524597167969
            im_multiplicator => "0010000110010011",
            data_re_out => mul_re_out(1835),
            data_im_out => mul_im_out(1835)
        );

 
    UMUL_1836 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1836),
            data_im_in => first_stage_im_out(1836),
            re_multiplicator => "1100110010011000", --- -0.80322265625 + j0.595703125
            im_multiplicator => "0010011000100000",
            data_re_out => mul_re_out(1836),
            data_im_out => mul_im_out(1836)
        );

 
    UMUL_1837 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1837),
            data_im_in => first_stage_im_out(1837),
            re_multiplicator => "1101000000001110", --- -0.749145507812 + j0.662414550781
            im_multiplicator => "0010101001100101",
            data_re_out => mul_re_out(1837),
            data_im_out => mul_im_out(1837)
        );

 
    UMUL_1838 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1838),
            data_im_in => first_stage_im_out(1838),
            re_multiplicator => "1101001111011111", --- -0.689514160156 + j0.724243164062
            im_multiplicator => "0010111001011010",
            data_re_out => mul_re_out(1838),
            data_im_out => mul_im_out(1838)
        );

 
    UMUL_1839 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1839),
            data_im_in => first_stage_im_out(1839),
            re_multiplicator => "1101100000000010", --- -0.624877929688 + j0.78076171875
            im_multiplicator => "0011000111111000",
            data_re_out => mul_re_out(1839),
            data_im_out => mul_im_out(1839)
        );

 
    UMUL_1840 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1840),
            data_im_in => first_stage_im_out(1840),
            re_multiplicator => "1101110001110010", --- -0.555541992188 + j0.831481933594
            im_multiplicator => "0011010100110111",
            data_re_out => mul_re_out(1840),
            data_im_out => mul_im_out(1840)
        );

 
    UMUL_1841 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1841),
            data_im_in => first_stage_im_out(1841),
            re_multiplicator => "1110000100100100", --- -0.482177734375 + j0.876098632812
            im_multiplicator => "0011100000010010",
            data_re_out => mul_re_out(1841),
            data_im_out => mul_im_out(1841)
        );

 
    UMUL_1842 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1842),
            data_im_in => first_stage_im_out(1842),
            re_multiplicator => "1110011000010001", --- -0.405212402344 + j0.914184570312
            im_multiplicator => "0011101010000010",
            data_re_out => mul_re_out(1842),
            data_im_out => mul_im_out(1842)
        );

 
    UMUL_1843 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1843),
            data_im_in => first_stage_im_out(1843),
            re_multiplicator => "1110101100101110", --- -0.325317382812 + j0.945617675781
            im_multiplicator => "0011110010000101",
            data_re_out => mul_re_out(1843),
            data_im_out => mul_im_out(1843)
        );

 
    UMUL_1844 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1844),
            data_im_in => first_stage_im_out(1844),
            re_multiplicator => "1111000001110011", --- -0.242980957031 + j0.970031738281
            im_multiplicator => "0011111000010101",
            data_re_out => mul_re_out(1844),
            data_im_out => mul_im_out(1844)
        );

 
    UMUL_1845 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1845),
            data_im_in => first_stage_im_out(1845),
            re_multiplicator => "1111010111010101", --- -0.158874511719 + j0.9873046875
            im_multiplicator => "0011111100110000",
            data_re_out => mul_re_out(1845),
            data_im_out => mul_im_out(1845)
        );

 
    UMUL_1846 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1846),
            data_im_in => first_stage_im_out(1846),
            re_multiplicator => "1111101101001011", --- -0.0735473632812 + j0.997314453125
            im_multiplicator => "0011111111010100",
            data_re_out => mul_re_out(1846),
            data_im_out => mul_im_out(1846)
        );

 
    UMUL_1847 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1847),
            data_im_in => first_stage_im_out(1847),
            re_multiplicator => "0000000011001001", --- 0.0122680664062 + j0.999938964844
            im_multiplicator => "0011111111111111",
            data_re_out => mul_re_out(1847),
            data_im_out => mul_im_out(1847)
        );

 
    UMUL_1848 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1848),
            data_im_in => first_stage_im_out(1848),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j0.995178222656
            im_multiplicator => "0011111110110001",
            data_re_out => mul_re_out(1848),
            data_im_out => mul_im_out(1848)
        );

 
    UMUL_1849 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1849),
            data_im_in => first_stage_im_out(1849),
            re_multiplicator => "0000101110110111", --- 0.183044433594 + j0.983093261719
            im_multiplicator => "0011111011101011",
            data_re_out => mul_re_out(1849),
            data_im_out => mul_im_out(1849)
        );

 
    UMUL_1850 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1850),
            data_im_in => first_stage_im_out(1850),
            re_multiplicator => "0001000100010010", --- 0.266723632812 + j0.963806152344
            im_multiplicator => "0011110110101111",
            data_re_out => mul_re_out(1850),
            data_im_out => mul_im_out(1850)
        );

 
    UMUL_1851 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1851),
            data_im_in => first_stage_im_out(1851),
            re_multiplicator => "0001011001001100", --- 0.348388671875 + j0.937316894531
            im_multiplicator => "0011101111111101",
            data_re_out => mul_re_out(1851),
            data_im_out => mul_im_out(1851)
        );

 
    UMUL_1852 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1852),
            data_im_in => first_stage_im_out(1852),
            re_multiplicator => "0001101101011101", --- 0.427551269531 + j0.903991699219
            im_multiplicator => "0011100111011011",
            data_re_out => mul_re_out(1852),
            data_im_out => mul_im_out(1852)
        );

 
    UMUL_1853 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1853),
            data_im_in => first_stage_im_out(1853),
            re_multiplicator => "0010000000111010", --- 0.503540039062 + j0.863952636719
            im_multiplicator => "0011011101001011",
            data_re_out => mul_re_out(1853),
            data_im_out => mul_im_out(1853)
        );

 
    UMUL_1854 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1854),
            data_im_in => first_stage_im_out(1854),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j0.817565917969
            im_multiplicator => "0011010001010011",
            data_re_out => mul_re_out(1854),
            data_im_out => mul_im_out(1854)
        );

 
    UMUL_1855 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1855),
            data_im_in => first_stage_im_out(1855),
            re_multiplicator => "0010100100110101", --- 0.643859863281 + j0.765197753906
            im_multiplicator => "0011000011111001",
            data_re_out => mul_re_out(1855),
            data_im_out => mul_im_out(1855)
        );

 
    UMUL_1856 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1856),
            data_im_in => first_stage_im_out(1856),
            data_re_out => mul_re_out(1856),
            data_im_out => mul_im_out(1856)
        );

 
    UMUL_1857 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1857),
            data_im_in => first_stage_im_out(1857),
            re_multiplicator => "0011111110111111", --- 0.996032714844 + j-0.0888671875
            im_multiplicator => "1111101001010000",
            data_re_out => mul_re_out(1857),
            data_im_out => mul_im_out(1857)
        );

 
    UMUL_1858 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1858),
            data_im_in => first_stage_im_out(1858),
            re_multiplicator => "0011111011111101", --- 0.984191894531 + j-0.177001953125
            im_multiplicator => "1111010010101100",
            data_re_out => mul_re_out(1858),
            data_im_out => mul_im_out(1858)
        );

 
    UMUL_1859 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1859),
            data_im_in => first_stage_im_out(1859),
            re_multiplicator => "0011110110111100", --- 0.964599609375 + j-0.263732910156
            im_multiplicator => "1110111100011111",
            data_re_out => mul_re_out(1859),
            data_im_out => mul_im_out(1859)
        );

 
    UMUL_1860 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1860),
            data_im_in => first_stage_im_out(1860),
            re_multiplicator => "0011101111111101", --- 0.937316894531 + j-0.348388671875
            im_multiplicator => "1110100110110100",
            data_re_out => mul_re_out(1860),
            data_im_out => mul_im_out(1860)
        );

 
    UMUL_1861 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1861),
            data_im_in => first_stage_im_out(1861),
            re_multiplicator => "0011100111000101", --- 0.902648925781 + j-0.430297851562
            im_multiplicator => "1110010001110110",
            data_re_out => mul_re_out(1861),
            data_im_out => mul_im_out(1861)
        );

 
    UMUL_1862 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1862),
            data_im_in => first_stage_im_out(1862),
            re_multiplicator => "0011011100011000", --- 0.86083984375 + j-0.508850097656
            im_multiplicator => "1101111101101111",
            data_re_out => mul_re_out(1862),
            data_im_out => mul_im_out(1862)
        );

 
    UMUL_1863 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1863),
            data_im_in => first_stage_im_out(1863),
            re_multiplicator => "0011001111111100", --- 0.812255859375 + j-0.583312988281
            im_multiplicator => "1101101010101011",
            data_re_out => mul_re_out(1863),
            data_im_out => mul_im_out(1863)
        );

 
    UMUL_1864 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1864),
            data_im_in => first_stage_im_out(1864),
            re_multiplicator => "0011000001110110", --- 0.757202148438 + j-0.653198242188
            im_multiplicator => "1101011000110010",
            data_re_out => mul_re_out(1864),
            data_im_out => mul_im_out(1864)
        );

 
    UMUL_1865 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1865),
            data_im_in => first_stage_im_out(1865),
            re_multiplicator => "0010110010001110", --- 0.696166992188 + j-0.717895507812
            im_multiplicator => "1101001000001110",
            data_re_out => mul_re_out(1865),
            data_im_out => mul_im_out(1865)
        );

 
    UMUL_1866 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1866),
            data_im_in => first_stage_im_out(1866),
            re_multiplicator => "0010100001001100", --- 0.629638671875 + j-0.776916503906
            im_multiplicator => "1100111001000111",
            data_re_out => mul_re_out(1866),
            data_im_out => mul_im_out(1866)
        );

 
    UMUL_1867 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1867),
            data_im_in => first_stage_im_out(1867),
            re_multiplicator => "0010001110111000", --- 0.55810546875 + j-0.829772949219
            im_multiplicator => "1100101011100101",
            data_re_out => mul_re_out(1867),
            data_im_out => mul_im_out(1867)
        );

 
    UMUL_1868 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1868),
            data_im_in => first_stage_im_out(1868),
            re_multiplicator => "0001111011011100", --- 0.482177734375 + j-0.876098632812
            im_multiplicator => "1100011111101110",
            data_re_out => mul_re_out(1868),
            data_im_out => mul_im_out(1868)
        );

 
    UMUL_1869 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1869),
            data_im_in => first_stage_im_out(1869),
            re_multiplicator => "0001100111000001", --- 0.402404785156 + j-0.915466308594
            im_multiplicator => "1100010101101001",
            data_re_out => mul_re_out(1869),
            data_im_out => mul_im_out(1869)
        );

 
    UMUL_1870 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1870),
            data_im_in => first_stage_im_out(1870),
            re_multiplicator => "0001010001110011", --- 0.319519042969 + j-0.947570800781
            im_multiplicator => "1100001101011011",
            data_re_out => mul_re_out(1870),
            data_im_out => mul_im_out(1870)
        );

 
    UMUL_1871 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1871),
            data_im_in => first_stage_im_out(1871),
            re_multiplicator => "0000111011111011", --- 0.234069824219 + j-0.972229003906
            im_multiplicator => "1100000111000111",
            data_re_out => mul_re_out(1871),
            data_im_out => mul_im_out(1871)
        );

 
    UMUL_1872 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1872),
            data_im_in => first_stage_im_out(1872),
            re_multiplicator => "0000100101100100", --- 0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(1872),
            data_im_out => mul_im_out(1872)
        );

 
    UMUL_1873 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1873),
            data_im_in => first_stage_im_out(1873),
            re_multiplicator => "0000001110111011", --- 0.0582885742188 + j-0.998291015625
            im_multiplicator => "1100000000011100",
            data_re_out => mul_re_out(1873),
            data_im_out => mul_im_out(1873)
        );

 
    UMUL_1874 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1874),
            data_im_in => first_stage_im_out(1874),
            re_multiplicator => "1111111000001001", --- -0.0307006835938 + j-0.99951171875
            im_multiplicator => "1100000000001000",
            data_re_out => mul_re_out(1874),
            data_im_out => mul_im_out(1874)
        );

 
    UMUL_1875 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1875),
            data_im_in => first_stage_im_out(1875),
            re_multiplicator => "1111100001011100", --- -0.119384765625 + j-0.992858886719
            im_multiplicator => "1100000001110101",
            data_re_out => mul_re_out(1875),
            data_im_out => mul_im_out(1875)
        );

 
    UMUL_1876 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1876),
            data_im_in => first_stage_im_out(1876),
            re_multiplicator => "1111001010111111", --- -0.207092285156 + j-0.978332519531
            im_multiplicator => "1100000101100011",
            data_re_out => mul_re_out(1876),
            data_im_out => mul_im_out(1876)
        );

 
    UMUL_1877 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1877),
            data_im_in => first_stage_im_out(1877),
            re_multiplicator => "1110110100111100", --- -0.293212890625 + j-0.9560546875
            im_multiplicator => "1100001011010000",
            data_re_out => mul_re_out(1877),
            data_im_out => mul_im_out(1877)
        );

 
    UMUL_1878 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1878),
            data_im_in => first_stage_im_out(1878),
            re_multiplicator => "1110011111011111", --- -0.377014160156 + j-0.926208496094
            im_multiplicator => "1100010010111001",
            data_re_out => mul_re_out(1878),
            data_im_out => mul_im_out(1878)
        );

 
    UMUL_1879 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1879),
            data_im_in => first_stage_im_out(1879),
            re_multiplicator => "1110001010110011", --- -0.457824707031 + j-0.889038085938
            im_multiplicator => "1100011100011010",
            data_re_out => mul_re_out(1879),
            data_im_out => mul_im_out(1879)
        );

 
    UMUL_1880 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1880),
            data_im_in => first_stage_im_out(1880),
            re_multiplicator => "1101110111000011", --- -0.534973144531 + j-0.844848632812
            im_multiplicator => "1100100111101110",
            data_re_out => mul_re_out(1880),
            data_im_out => mul_im_out(1880)
        );

 
    UMUL_1881 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1881),
            data_im_in => first_stage_im_out(1881),
            re_multiplicator => "1101100100010111", --- -0.607971191406 + j-0.7939453125
            im_multiplicator => "1100110100110000",
            data_re_out => mul_re_out(1881),
            data_im_out => mul_im_out(1881)
        );

 
    UMUL_1882 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1882),
            data_im_in => first_stage_im_out(1882),
            re_multiplicator => "1101010010111011", --- -0.676086425781 + j-0.73681640625
            im_multiplicator => "1101000011011000",
            data_re_out => mul_re_out(1882),
            data_im_out => mul_im_out(1882)
        );

 
    UMUL_1883 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1883),
            data_im_in => first_stage_im_out(1883),
            re_multiplicator => "1101000010110110", --- -0.738891601562 + j-0.673828125
            im_multiplicator => "1101010011100000",
            data_re_out => mul_re_out(1883),
            data_im_out => mul_im_out(1883)
        );

 
    UMUL_1884 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1884),
            data_im_in => first_stage_im_out(1884),
            re_multiplicator => "1100110100010001", --- -0.795837402344 + j-0.605529785156
            im_multiplicator => "1101100100111111",
            data_re_out => mul_re_out(1884),
            data_im_out => mul_im_out(1884)
        );

 
    UMUL_1885 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1885),
            data_im_in => first_stage_im_out(1885),
            re_multiplicator => "1100100111010011", --- -0.846496582031 + j-0.532409667969
            im_multiplicator => "1101110111101101",
            data_re_out => mul_re_out(1885),
            data_im_out => mul_im_out(1885)
        );

 
    UMUL_1886 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1886),
            data_im_in => first_stage_im_out(1886),
            re_multiplicator => "1100011100000011", --- -0.890441894531 + j-0.455078125
            im_multiplicator => "1110001011100000",
            data_re_out => mul_re_out(1886),
            data_im_out => mul_im_out(1886)
        );

 
    UMUL_1887 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1887),
            data_im_in => first_stage_im_out(1887),
            re_multiplicator => "1100010010100110", --- -0.927368164062 + j-0.374145507812
            im_multiplicator => "1110100000001110",
            data_re_out => mul_re_out(1887),
            data_im_out => mul_im_out(1887)
        );

 
    UMUL_1888 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1888),
            data_im_in => first_stage_im_out(1888),
            re_multiplicator => "1100001011000001", --- -0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(1888),
            data_im_out => mul_im_out(1888)
        );

 
    UMUL_1889 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1889),
            data_im_in => first_stage_im_out(1889),
            re_multiplicator => "1100000101011001", --- -0.978942871094 + j-0.2041015625
            im_multiplicator => "1111001011110000",
            data_re_out => mul_re_out(1889),
            data_im_out => mul_im_out(1889)
        );

 
    UMUL_1890 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1890),
            data_im_in => first_stage_im_out(1890),
            re_multiplicator => "1100000001101111", --- -0.993225097656 + j-0.116333007812
            im_multiplicator => "1111100010001110",
            data_re_out => mul_re_out(1890),
            data_im_out => mul_im_out(1890)
        );

 
    UMUL_1891 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1891),
            data_im_in => first_stage_im_out(1891),
            re_multiplicator => "1100000000000110", --- -0.999633789062 + j-0.027587890625
            im_multiplicator => "1111111000111100",
            data_re_out => mul_re_out(1891),
            data_im_out => mul_im_out(1891)
        );

 
    UMUL_1892 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1892),
            data_im_in => first_stage_im_out(1892),
            re_multiplicator => "1100000000011111", --- -0.998107910156 + j0.0613403320312
            im_multiplicator => "0000001111101101",
            data_re_out => mul_re_out(1892),
            data_im_out => mul_im_out(1892)
        );

 
    UMUL_1893 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1893),
            data_im_in => first_stage_im_out(1893),
            re_multiplicator => "1100000010111001", --- -0.988708496094 + j0.149780273438
            im_multiplicator => "0000100110010110",
            data_re_out => mul_re_out(1893),
            data_im_out => mul_im_out(1893)
        );

 
    UMUL_1894 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1894),
            data_im_in => first_stage_im_out(1894),
            re_multiplicator => "1100000111010011", --- -0.971496582031 + j0.236999511719
            im_multiplicator => "0000111100101011",
            data_re_out => mul_re_out(1894),
            data_im_out => mul_im_out(1894)
        );

 
    UMUL_1895 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1895),
            data_im_in => first_stage_im_out(1895),
            re_multiplicator => "1100001101101011", --- -0.946594238281 + j0.322387695312
            im_multiplicator => "0001010010100010",
            data_re_out => mul_re_out(1895),
            data_im_out => mul_im_out(1895)
        );

 
    UMUL_1896 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1896),
            data_im_in => first_stage_im_out(1896),
            re_multiplicator => "1100010101111110", --- -0.914184570312 + j0.405212402344
            im_multiplicator => "0001100111101111",
            data_re_out => mul_re_out(1896),
            data_im_out => mul_im_out(1896)
        );

 
    UMUL_1897 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1897),
            data_im_in => first_stage_im_out(1897),
            re_multiplicator => "1100100000000111", --- -0.874572753906 + j0.48486328125
            im_multiplicator => "0001111100001000",
            data_re_out => mul_re_out(1897),
            data_im_out => mul_im_out(1897)
        );

 
    UMUL_1898 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1898),
            data_im_in => first_stage_im_out(1898),
            re_multiplicator => "1100101100000001", --- -0.828063964844 + j0.560668945312
            im_multiplicator => "0010001111100010",
            data_re_out => mul_re_out(1898),
            data_im_out => mul_im_out(1898)
        );

 
    UMUL_1899 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1899),
            data_im_in => first_stage_im_out(1899),
            re_multiplicator => "1100111001100111", --- -0.774963378906 + j0.632019042969
            im_multiplicator => "0010100001110011",
            data_re_out => mul_re_out(1899),
            data_im_out => mul_im_out(1899)
        );

 
    UMUL_1900 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1900),
            data_im_in => first_stage_im_out(1900),
            re_multiplicator => "1101001000110001", --- -0.715759277344 + j0.698364257812
            im_multiplicator => "0010110010110010",
            data_re_out => mul_re_out(1900),
            data_im_out => mul_im_out(1900)
        );

 
    UMUL_1901 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1901),
            data_im_in => first_stage_im_out(1901),
            re_multiplicator => "1101011001011001", --- -0.650817871094 + j0.759216308594
            im_multiplicator => "0011000010010111",
            data_re_out => mul_re_out(1901),
            data_im_out => mul_im_out(1901)
        );

 
    UMUL_1902 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1902),
            data_im_in => first_stage_im_out(1902),
            re_multiplicator => "1101101011010100", --- -0.580810546875 + j0.814025878906
            im_multiplicator => "0011010000011001",
            data_re_out => mul_re_out(1902),
            data_im_out => mul_im_out(1902)
        );

 
    UMUL_1903 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1903),
            data_im_in => first_stage_im_out(1903),
            re_multiplicator => "1101111110011011", --- -0.506164550781 + j0.862426757812
            im_multiplicator => "0011011100110010",
            data_re_out => mul_re_out(1903),
            data_im_out => mul_im_out(1903)
        );

 
    UMUL_1904 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1904),
            data_im_in => first_stage_im_out(1904),
            re_multiplicator => "1110010010100011", --- -0.427551269531 + j0.903991699219
            im_multiplicator => "0011100111011011",
            data_re_out => mul_re_out(1904),
            data_im_out => mul_im_out(1904)
        );

 
    UMUL_1905 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1905),
            data_im_in => first_stage_im_out(1905),
            re_multiplicator => "1110100111100011", --- -0.345520019531 + j0.938415527344
            im_multiplicator => "0011110000001111",
            data_re_out => mul_re_out(1905),
            data_im_out => mul_im_out(1905)
        );

 
    UMUL_1906 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1906),
            data_im_in => first_stage_im_out(1906),
            re_multiplicator => "1110111101001111", --- -0.260803222656 + j0.965393066406
            im_multiplicator => "0011110111001001",
            data_re_out => mul_re_out(1906),
            data_im_out => mul_im_out(1906)
        );

 
    UMUL_1907 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1907),
            data_im_in => first_stage_im_out(1907),
            re_multiplicator => "1111010011011101", --- -0.174011230469 + j0.984741210938
            im_multiplicator => "0011111100000110",
            data_re_out => mul_re_out(1907),
            data_im_out => mul_im_out(1907)
        );

 
    UMUL_1908 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1908),
            data_im_in => first_stage_im_out(1908),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j0.996337890625
            im_multiplicator => "0011111111000100",
            data_re_out => mul_re_out(1908),
            data_im_out => mul_im_out(1908)
        );

 
    UMUL_1909 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1909),
            data_im_in => first_stage_im_out(1909),
            re_multiplicator => "0000000000110010", --- 0.0030517578125 + j1.0
            im_multiplicator => "0100000000000000",
            data_re_out => mul_re_out(1909),
            data_im_out => mul_im_out(1909)
        );

 
    UMUL_1910 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1910),
            data_im_in => first_stage_im_out(1910),
            re_multiplicator => "0000010111100010", --- 0.0919189453125 + j0.995788574219
            im_multiplicator => "0011111110111011",
            data_re_out => mul_re_out(1910),
            data_im_out => mul_im_out(1910)
        );

 
    UMUL_1911 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1911),
            data_im_in => first_stage_im_out(1911),
            re_multiplicator => "0000101110000101", --- 0.179992675781 + j0.983642578125
            im_multiplicator => "0011111011110100",
            data_re_out => mul_re_out(1911),
            data_im_out => mul_im_out(1911)
        );

 
    UMUL_1912 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1912),
            data_im_in => first_stage_im_out(1912),
            re_multiplicator => "0001000100010010", --- 0.266723632812 + j0.963806152344
            im_multiplicator => "0011110110101111",
            data_re_out => mul_re_out(1912),
            data_im_out => mul_im_out(1912)
        );

 
    UMUL_1913 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1913),
            data_im_in => first_stage_im_out(1913),
            re_multiplicator => "0001011001111100", --- 0.351318359375 + j0.936279296875
            im_multiplicator => "0011101111101100",
            data_re_out => mul_re_out(1913),
            data_im_out => mul_im_out(1913)
        );

 
    UMUL_1914 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1914),
            data_im_in => first_stage_im_out(1914),
            re_multiplicator => "0001101110111000", --- 0.43310546875 + j0.9013671875
            im_multiplicator => "0011100110110000",
            data_re_out => mul_re_out(1914),
            data_im_out => mul_im_out(1914)
        );

 
    UMUL_1915 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1915),
            data_im_in => first_stage_im_out(1915),
            re_multiplicator => "0010000010111100", --- 0.511474609375 + j0.859313964844
            im_multiplicator => "0011011011111111",
            data_re_out => mul_re_out(1915),
            data_im_out => mul_im_out(1915)
        );

 
    UMUL_1916 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1916),
            data_im_in => first_stage_im_out(1916),
            re_multiplicator => "0010010101111110", --- 0.585815429688 + j0.810485839844
            im_multiplicator => "0011001111011111",
            data_re_out => mul_re_out(1916),
            data_im_out => mul_im_out(1916)
        );

 
    UMUL_1917 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1917),
            data_im_in => first_stage_im_out(1917),
            re_multiplicator => "0010100111110100", --- 0.655517578125 + j0.755187988281
            im_multiplicator => "0011000001010101",
            data_re_out => mul_re_out(1917),
            data_im_out => mul_im_out(1917)
        );

 
    UMUL_1918 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1918),
            data_im_in => first_stage_im_out(1918),
            re_multiplicator => "0010111000010101", --- 0.720031738281 + j0.693969726562
            im_multiplicator => "0010110001101010",
            data_re_out => mul_re_out(1918),
            data_im_out => mul_im_out(1918)
        );

 
    UMUL_1919 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1919),
            data_im_in => first_stage_im_out(1919),
            re_multiplicator => "0011000111011000", --- 0.77880859375 + j0.627258300781
            im_multiplicator => "0010100000100101",
            data_re_out => mul_re_out(1919),
            data_im_out => mul_im_out(1919)
        );

 
    UMUL_1920 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1920),
            data_im_in => first_stage_im_out(1920),
            data_re_out => mul_re_out(1920),
            data_im_out => mul_im_out(1920)
        );

 
    UMUL_1921 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1921),
            data_im_in => first_stage_im_out(1921),
            re_multiplicator => "0011111110111011", --- 0.995788574219 + j-0.0919189453125
            im_multiplicator => "1111101000011110",
            data_re_out => mul_re_out(1921),
            data_im_out => mul_im_out(1921)
        );

 
    UMUL_1922 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1922),
            data_im_in => first_stage_im_out(1922),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(1922),
            data_im_out => mul_im_out(1922)
        );

 
    UMUL_1923 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1923),
            data_im_in => first_stage_im_out(1923),
            re_multiplicator => "0011110110010011", --- 0.962097167969 + j-0.272644042969
            im_multiplicator => "1110111010001101",
            data_re_out => mul_re_out(1923),
            data_im_out => mul_im_out(1923)
        );

 
    UMUL_1924 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1924),
            data_im_in => first_stage_im_out(1924),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(1924),
            data_im_out => mul_im_out(1924)
        );

 
    UMUL_1925 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1925),
            data_im_in => first_stage_im_out(1925),
            re_multiplicator => "0011100101011000", --- 0.89599609375 + j-0.444091796875
            im_multiplicator => "1110001110010100",
            data_re_out => mul_re_out(1925),
            data_im_out => mul_im_out(1925)
        );

 
    UMUL_1926 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1926),
            data_im_in => first_stage_im_out(1926),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(1926),
            data_im_out => mul_im_out(1926)
        );

 
    UMUL_1927 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1927),
            data_im_in => first_stage_im_out(1927),
            re_multiplicator => "0011001100101100", --- 0.799560546875 + j-0.600646972656
            im_multiplicator => "1101100110001111",
            data_re_out => mul_re_out(1927),
            data_im_out => mul_im_out(1927)
        );

 
    UMUL_1928 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1928),
            data_im_in => first_stage_im_out(1928),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(1928),
            data_im_out => mul_im_out(1928)
        );

 
    UMUL_1929 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1929),
            data_im_in => first_stage_im_out(1929),
            re_multiplicator => "0010101101000101", --- 0.676086425781 + j-0.73681640625
            im_multiplicator => "1101000011011000",
            data_re_out => mul_re_out(1929),
            data_im_out => mul_im_out(1929)
        );

 
    UMUL_1930 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1930),
            data_im_in => first_stage_im_out(1930),
            re_multiplicator => "0010011011000001", --- 0.605529785156 + j-0.795837402344
            im_multiplicator => "1100110100010001",
            data_re_out => mul_re_out(1930),
            data_im_out => mul_im_out(1930)
        );

 
    UMUL_1931 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1931),
            data_im_in => first_stage_im_out(1931),
            re_multiplicator => "0010000111101000", --- 0.52978515625 + j-0.84814453125
            im_multiplicator => "1100100110111000",
            data_re_out => mul_re_out(1931),
            data_im_out => mul_im_out(1931)
        );

 
    UMUL_1932 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1932),
            data_im_in => first_stage_im_out(1932),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(1932),
            data_im_out => mul_im_out(1932)
        );

 
    UMUL_1933 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1933),
            data_im_in => first_stage_im_out(1933),
            re_multiplicator => "0001011101100110", --- 0.365600585938 + j-0.930786132812
            im_multiplicator => "1100010001101110",
            data_re_out => mul_re_out(1933),
            data_im_out => mul_im_out(1933)
        );

 
    UMUL_1934 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1934),
            data_im_in => first_stage_im_out(1934),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(1934),
            data_im_out => mul_im_out(1934)
        );

 
    UMUL_1935 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1935),
            data_im_in => first_stage_im_out(1935),
            re_multiplicator => "0000110000011010", --- 0.189086914062 + j-0.98193359375
            im_multiplicator => "1100000100101000",
            data_re_out => mul_re_out(1935),
            data_im_out => mul_im_out(1935)
        );

 
    UMUL_1936 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1936),
            data_im_in => first_stage_im_out(1936),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(1936),
            data_im_out => mul_im_out(1936)
        );

 
    UMUL_1937 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1937),
            data_im_in => first_stage_im_out(1937),
            re_multiplicator => "0000000001100101", --- 0.00616455078125 + j-1.0
            im_multiplicator => "1100000000000000",
            data_re_out => mul_re_out(1937),
            data_im_out => mul_im_out(1937)
        );

 
    UMUL_1938 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1938),
            data_im_in => first_stage_im_out(1938),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(1938),
            data_im_out => mul_im_out(1938)
        );

 
    UMUL_1939 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1939),
            data_im_in => first_stage_im_out(1939),
            re_multiplicator => "1111010010101100", --- -0.177001953125 + j-0.984191894531
            im_multiplicator => "1100000100000011",
            data_re_out => mul_re_out(1939),
            data_im_out => mul_im_out(1939)
        );

 
    UMUL_1940 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1940),
            data_im_in => first_stage_im_out(1940),
            re_multiplicator => "1110111011101110", --- -0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(1940),
            data_im_out => mul_im_out(1940)
        );

 
    UMUL_1941 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1941),
            data_im_in => first_stage_im_out(1941),
            re_multiplicator => "1110100101010101", --- -0.354187011719 + j-0.935180664062
            im_multiplicator => "1100010000100110",
            data_re_out => mul_re_out(1941),
            data_im_out => mul_im_out(1941)
        );

 
    UMUL_1942 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1942),
            data_im_in => first_stage_im_out(1942),
            re_multiplicator => "1110001111101110", --- -0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(1942),
            data_im_out => mul_im_out(1942)
        );

 
    UMUL_1943 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1943),
            data_im_in => first_stage_im_out(1943),
            re_multiplicator => "1101111011000011", --- -0.519348144531 + j-0.854553222656
            im_multiplicator => "1100100101001111",
            data_re_out => mul_re_out(1943),
            data_im_out => mul_im_out(1943)
        );

 
    UMUL_1944 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1944),
            data_im_in => first_stage_im_out(1944),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(1944),
            data_im_out => mul_im_out(1944)
        );

 
    UMUL_1945 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1945),
            data_im_in => first_stage_im_out(1945),
            re_multiplicator => "1101010101010000", --- -0.6669921875 + j-0.745056152344
            im_multiplicator => "1101000001010001",
            data_re_out => mul_re_out(1945),
            data_im_out => mul_im_out(1945)
        );

 
    UMUL_1946 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1946),
            data_im_in => first_stage_im_out(1946),
            re_multiplicator => "1101000100011100", --- -0.732666015625 + j-0.680603027344
            im_multiplicator => "1101010001110001",
            data_re_out => mul_re_out(1946),
            data_im_out => mul_im_out(1946)
        );

 
    UMUL_1947 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1947),
            data_im_in => first_stage_im_out(1947),
            re_multiplicator => "1100110101001110", --- -0.792114257812 + j-0.610412597656
            im_multiplicator => "1101100011101111",
            data_re_out => mul_re_out(1947),
            data_im_out => mul_im_out(1947)
        );

 
    UMUL_1948 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1948),
            data_im_in => first_stage_im_out(1948),
            re_multiplicator => "1100100111101110", --- -0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(1948),
            data_im_out => mul_im_out(1948)
        );

 
    UMUL_1949 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1949),
            data_im_in => first_stage_im_out(1949),
            re_multiplicator => "1100011100000011", --- -0.890441894531 + j-0.455078125
            im_multiplicator => "1110001011100000",
            data_re_out => mul_re_out(1949),
            data_im_out => mul_im_out(1949)
        );

 
    UMUL_1950 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1950),
            data_im_in => first_stage_im_out(1950),
            re_multiplicator => "1100010010010011", --- -0.928527832031 + j-0.371337890625
            im_multiplicator => "1110100000111100",
            data_re_out => mul_re_out(1950),
            data_im_out => mul_im_out(1950)
        );

 
    UMUL_1951 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1951),
            data_im_in => first_stage_im_out(1951),
            re_multiplicator => "1100001010100101", --- -0.958679199219 + j-0.284423828125
            im_multiplicator => "1110110111001100",
            data_re_out => mul_re_out(1951),
            data_im_out => mul_im_out(1951)
        );

 
    UMUL_1952 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1952),
            data_im_in => first_stage_im_out(1952),
            re_multiplicator => "1100000100111011", --- -0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(1952),
            data_im_out => mul_im_out(1952)
        );

 
    UMUL_1953 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1953),
            data_im_in => first_stage_im_out(1953),
            re_multiplicator => "1100000001011001", --- -0.994567871094 + j-0.104125976562
            im_multiplicator => "1111100101010110",
            data_re_out => mul_re_out(1953),
            data_im_out => mul_im_out(1953)
        );

 
    UMUL_1954 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1954),
            data_im_in => first_stage_im_out(1954),
            re_multiplicator => "1100000000000001", --- -0.999938964844 + j-0.0122680664062
            im_multiplicator => "1111111100110111",
            data_re_out => mul_re_out(1954),
            data_im_out => mul_im_out(1954)
        );

 
    UMUL_1955 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1955),
            data_im_in => first_stage_im_out(1955),
            re_multiplicator => "1100000000110100", --- -0.996826171875 + j0.0797119140625
            im_multiplicator => "0000010100011010",
            data_re_out => mul_re_out(1955),
            data_im_out => mul_im_out(1955)
        );

 
    UMUL_1956 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1956),
            data_im_in => first_stage_im_out(1956),
            re_multiplicator => "1100000011110001", --- -0.985290527344 + j0.170959472656
            im_multiplicator => "0000101011110001",
            data_re_out => mul_re_out(1956),
            data_im_out => mul_im_out(1956)
        );

 
    UMUL_1957 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1957),
            data_im_in => first_stage_im_out(1957),
            re_multiplicator => "1100001000110111", --- -0.965393066406 + j0.260803222656
            im_multiplicator => "0001000010110001",
            data_re_out => mul_re_out(1957),
            data_im_out => mul_im_out(1957)
        );

 
    UMUL_1958 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1958),
            data_im_in => first_stage_im_out(1958),
            re_multiplicator => "1100010000000011", --- -0.937316894531 + j0.348388671875
            im_multiplicator => "0001011001001100",
            data_re_out => mul_re_out(1958),
            data_im_out => mul_im_out(1958)
        );

 
    UMUL_1959 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1959),
            data_im_in => first_stage_im_out(1959),
            re_multiplicator => "1100011001010000", --- -0.9013671875 + j0.43310546875
            im_multiplicator => "0001101110111000",
            data_re_out => mul_re_out(1959),
            data_im_out => mul_im_out(1959)
        );

 
    UMUL_1960 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1960),
            data_im_in => first_stage_im_out(1960),
            re_multiplicator => "1100100100011011", --- -0.857727050781 + j0.514099121094
            im_multiplicator => "0010000011100111",
            data_re_out => mul_re_out(1960),
            data_im_out => mul_im_out(1960)
        );

 
    UMUL_1961 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1961),
            data_im_in => first_stage_im_out(1961),
            re_multiplicator => "1100110001011101", --- -0.806823730469 + j0.590759277344
            im_multiplicator => "0010010111001111",
            data_re_out => mul_re_out(1961),
            data_im_out => mul_im_out(1961)
        );

 
    UMUL_1962 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1962),
            data_im_in => first_stage_im_out(1962),
            re_multiplicator => "1101000000001110", --- -0.749145507812 + j0.662414550781
            im_multiplicator => "0010101001100101",
            data_re_out => mul_re_out(1962),
            data_im_out => mul_im_out(1962)
        );

 
    UMUL_1963 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1963),
            data_im_in => first_stage_im_out(1963),
            re_multiplicator => "1101010000101000", --- -0.68505859375 + j0.728454589844
            im_multiplicator => "0010111010011111",
            data_re_out => mul_re_out(1963),
            data_im_out => mul_im_out(1963)
        );

 
    UMUL_1964 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1964),
            data_im_in => first_stage_im_out(1964),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j0.788330078125
            im_multiplicator => "0011001001110100",
            data_re_out => mul_re_out(1964),
            data_im_out => mul_im_out(1964)
        );

 
    UMUL_1965 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1965),
            data_im_in => first_stage_im_out(1965),
            re_multiplicator => "1101110101101110", --- -0.540161132812 + j0.841552734375
            im_multiplicator => "0011010111011100",
            data_re_out => mul_re_out(1965),
            data_im_out => mul_im_out(1965)
        );

 
    UMUL_1966 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1966),
            data_im_in => first_stage_im_out(1966),
            re_multiplicator => "1110001010000111", --- -0.460510253906 + j0.887634277344
            im_multiplicator => "0011100011001111",
            data_re_out => mul_re_out(1966),
            data_im_out => mul_im_out(1966)
        );

 
    UMUL_1967 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1967),
            data_im_in => first_stage_im_out(1967),
            re_multiplicator => "1110011111011111", --- -0.377014160156 + j0.926208496094
            im_multiplicator => "0011101101000111",
            data_re_out => mul_re_out(1967),
            data_im_out => mul_im_out(1967)
        );

 
    UMUL_1968 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1968),
            data_im_in => first_stage_im_out(1968),
            re_multiplicator => "1110110101101100", --- -0.290283203125 + j0.956970214844
            im_multiplicator => "0011110100111111",
            data_re_out => mul_re_out(1968),
            data_im_out => mul_im_out(1968)
        );

 
    UMUL_1969 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1969),
            data_im_in => first_stage_im_out(1969),
            re_multiplicator => "1111001100100001", --- -0.201110839844 + j0.979553222656
            im_multiplicator => "0011111010110001",
            data_re_out => mul_re_out(1969),
            data_im_out => mul_im_out(1969)
        );

 
    UMUL_1970 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1970),
            data_im_in => first_stage_im_out(1970),
            re_multiplicator => "1111100011110010", --- -0.110229492188 + j0.993896484375
            im_multiplicator => "0011111110011100",
            data_re_out => mul_re_out(1970),
            data_im_out => mul_im_out(1970)
        );

 
    UMUL_1971 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1971),
            data_im_in => first_stage_im_out(1971),
            re_multiplicator => "1111111011010010", --- -0.0184326171875 + j0.999816894531
            im_multiplicator => "0011111111111101",
            data_re_out => mul_re_out(1971),
            data_im_out => mul_im_out(1971)
        );

 
    UMUL_1972 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1972),
            data_im_in => first_stage_im_out(1972),
            re_multiplicator => "0000010010110101", --- 0.0735473632812 + j0.997314453125
            im_multiplicator => "0011111111010100",
            data_re_out => mul_re_out(1972),
            data_im_out => mul_im_out(1972)
        );

 
    UMUL_1973 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1973),
            data_im_in => first_stage_im_out(1973),
            re_multiplicator => "0000101010001110", --- 0.164916992188 + j0.986328125
            im_multiplicator => "0011111100100000",
            data_re_out => mul_re_out(1973),
            data_im_out => mul_im_out(1973)
        );

 
    UMUL_1974 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1974),
            data_im_in => first_stage_im_out(1974),
            re_multiplicator => "0001000001010000", --- 0.2548828125 + j0.966979980469
            im_multiplicator => "0011110111100011",
            data_re_out => mul_re_out(1974),
            data_im_out => mul_im_out(1974)
        );

 
    UMUL_1975 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1975),
            data_im_in => first_stage_im_out(1975),
            re_multiplicator => "0001010111101110", --- 0.342651367188 + j0.939453125
            im_multiplicator => "0011110000100000",
            data_re_out => mul_re_out(1975),
            data_im_out => mul_im_out(1975)
        );

 
    UMUL_1976 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1976),
            data_im_in => first_stage_im_out(1976),
            re_multiplicator => "0001101101011101", --- 0.427551269531 + j0.903991699219
            im_multiplicator => "0011100111011011",
            data_re_out => mul_re_out(1976),
            data_im_out => mul_im_out(1976)
        );

 
    UMUL_1977 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1977),
            data_im_in => first_stage_im_out(1977),
            re_multiplicator => "0010000010010001", --- 0.508850097656 + j0.86083984375
            im_multiplicator => "0011011100011000",
            data_re_out => mul_re_out(1977),
            data_im_out => mul_im_out(1977)
        );

 
    UMUL_1978 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1978),
            data_im_in => first_stage_im_out(1978),
            re_multiplicator => "0010010101111110", --- 0.585815429688 + j0.810485839844
            im_multiplicator => "0011001111011111",
            data_re_out => mul_re_out(1978),
            data_im_out => mul_im_out(1978)
        );

 
    UMUL_1979 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1979),
            data_im_in => first_stage_im_out(1979),
            re_multiplicator => "0010101000011010", --- 0.657836914062 + j0.753173828125
            im_multiplicator => "0011000000110100",
            data_re_out => mul_re_out(1979),
            data_im_out => mul_im_out(1979)
        );

 
    UMUL_1980 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1980),
            data_im_in => first_stage_im_out(1980),
            re_multiplicator => "0010111001011010", --- 0.724243164062 + j0.689514160156
            im_multiplicator => "0010110000100001",
            data_re_out => mul_re_out(1980),
            data_im_out => mul_im_out(1980)
        );

 
    UMUL_1981 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1981),
            data_im_in => first_stage_im_out(1981),
            re_multiplicator => "0011001000110110", --- 0.784545898438 + j0.620056152344
            im_multiplicator => "0010011110101111",
            data_re_out => mul_re_out(1981),
            data_im_out => mul_im_out(1981)
        );

 
    UMUL_1982 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1982),
            data_im_in => first_stage_im_out(1982),
            re_multiplicator => "0011010110100101", --- 0.838195800781 + j0.545349121094
            im_multiplicator => "0010001011100111",
            data_re_out => mul_re_out(1982),
            data_im_out => mul_im_out(1982)
        );

 
    UMUL_1983 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1983),
            data_im_in => first_stage_im_out(1983),
            re_multiplicator => "0011100010100001", --- 0.884826660156 + j0.466003417969
            im_multiplicator => "0001110111010011",
            data_re_out => mul_re_out(1983),
            data_im_out => mul_im_out(1983)
        );

 
    UMUL_1984 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1984),
            data_im_in => first_stage_im_out(1984),
            data_re_out => mul_re_out(1984),
            data_im_out => mul_im_out(1984)
        );

 
    UMUL_1985 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1985),
            data_im_in => first_stage_im_out(1985),
            re_multiplicator => "0011111110110110", --- 0.995483398438 + j-0.094970703125
            im_multiplicator => "1111100111101100",
            data_re_out => mul_re_out(1985),
            data_im_out => mul_im_out(1985)
        );

 
    UMUL_1986 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1986),
            data_im_in => first_stage_im_out(1986),
            re_multiplicator => "0011111011011000", --- 0.98193359375 + j-0.189086914062
            im_multiplicator => "1111001111100110",
            data_re_out => mul_re_out(1986),
            data_im_out => mul_im_out(1986)
        );

 
    UMUL_1987 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1987),
            data_im_in => first_stage_im_out(1987),
            re_multiplicator => "0011110101101010", --- 0.959594726562 + j-0.281494140625
            im_multiplicator => "1110110111111100",
            data_re_out => mul_re_out(1987),
            data_im_out => mul_im_out(1987)
        );

 
    UMUL_1988 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1988),
            data_im_in => first_stage_im_out(1988),
            re_multiplicator => "0011101101101101", --- 0.928527832031 + j-0.371337890625
            im_multiplicator => "1110100000111100",
            data_re_out => mul_re_out(1988),
            data_im_out => mul_im_out(1988)
        );

 
    UMUL_1989 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1989),
            data_im_in => first_stage_im_out(1989),
            re_multiplicator => "0011100011100110", --- 0.889038085938 + j-0.457824707031
            im_multiplicator => "1110001010110011",
            data_re_out => mul_re_out(1989),
            data_im_out => mul_im_out(1989)
        );

 
    UMUL_1990 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1990),
            data_im_in => first_stage_im_out(1990),
            re_multiplicator => "0011010111011100", --- 0.841552734375 + j-0.540161132812
            im_multiplicator => "1101110101101110",
            data_re_out => mul_re_out(1990),
            data_im_out => mul_im_out(1990)
        );

 
    UMUL_1991 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1991),
            data_im_in => first_stage_im_out(1991),
            re_multiplicator => "0011001001010101", --- 0.786437988281 + j-0.61767578125
            im_multiplicator => "1101100001111000",
            data_re_out => mul_re_out(1991),
            data_im_out => mul_im_out(1991)
        );

 
    UMUL_1992 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1992),
            data_im_in => first_stage_im_out(1992),
            re_multiplicator => "0010111001011010", --- 0.724243164062 + j-0.689514160156
            im_multiplicator => "1101001111011111",
            data_re_out => mul_re_out(1992),
            data_im_out => mul_im_out(1992)
        );

 
    UMUL_1993 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1993),
            data_im_in => first_stage_im_out(1993),
            re_multiplicator => "0010100111110100", --- 0.655517578125 + j-0.755187988281
            im_multiplicator => "1100111110101011",
            data_re_out => mul_re_out(1993),
            data_im_out => mul_im_out(1993)
        );

 
    UMUL_1994 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1994),
            data_im_in => first_stage_im_out(1994),
            re_multiplicator => "0010010100101100", --- 0.580810546875 + j-0.814025878906
            im_multiplicator => "1100101111100111",
            data_re_out => mul_re_out(1994),
            data_im_out => mul_im_out(1994)
        );

 
    UMUL_1995 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1995),
            data_im_in => first_stage_im_out(1995),
            re_multiplicator => "0010000000001111", --- 0.500915527344 + j-0.865539550781
            im_multiplicator => "1100100010011011",
            data_re_out => mul_re_out(1995),
            data_im_out => mul_im_out(1995)
        );

 
    UMUL_1996 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1996),
            data_im_in => first_stage_im_out(1996),
            re_multiplicator => "0001101010100111", --- 0.416442871094 + j-0.9091796875
            im_multiplicator => "1100010111010000",
            data_re_out => mul_re_out(1996),
            data_im_out => mul_im_out(1996)
        );

 
    UMUL_1997 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1997),
            data_im_in => first_stage_im_out(1997),
            re_multiplicator => "0001010100000001", --- 0.328186035156 + j-0.944580078125
            im_multiplicator => "1100001110001100",
            data_re_out => mul_re_out(1997),
            data_im_out => mul_im_out(1997)
        );

 
    UMUL_1998 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1998),
            data_im_in => first_stage_im_out(1998),
            re_multiplicator => "0000111100101011", --- 0.236999511719 + j-0.971496582031
            im_multiplicator => "1100000111010011",
            data_re_out => mul_re_out(1998),
            data_im_out => mul_im_out(1998)
        );

 
    UMUL_1999 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1999),
            data_im_in => first_stage_im_out(1999),
            re_multiplicator => "0000100100110010", --- 0.143676757812 + j-0.989624023438
            im_multiplicator => "1100000010101010",
            data_re_out => mul_re_out(1999),
            data_im_out => mul_im_out(1999)
        );

 
    UMUL_2000 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2000),
            data_im_in => first_stage_im_out(2000),
            re_multiplicator => "0000001100100100", --- 0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(2000),
            data_im_out => mul_im_out(2000)
        );

 
    UMUL_2001 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2001),
            data_im_in => first_stage_im_out(2001),
            re_multiplicator => "1111110100001110", --- -0.0460205078125 + j-0.998962402344
            im_multiplicator => "1100000000010001",
            data_re_out => mul_re_out(2001),
            data_im_out => mul_im_out(2001)
        );

 
    UMUL_2002 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2002),
            data_im_in => first_stage_im_out(2002),
            re_multiplicator => "1111011011111111", --- -0.140686035156 + j-0.990051269531
            im_multiplicator => "1100000010100011",
            data_re_out => mul_re_out(2002),
            data_im_out => mul_im_out(2002)
        );

 
    UMUL_2003 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2003),
            data_im_in => first_stage_im_out(2003),
            re_multiplicator => "1111000100000101", --- -0.234069824219 + j-0.972229003906
            im_multiplicator => "1100000111000111",
            data_re_out => mul_re_out(2003),
            data_im_out => mul_im_out(2003)
        );

 
    UMUL_2004 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2004),
            data_im_in => first_stage_im_out(2004),
            re_multiplicator => "1110101100101110", --- -0.325317382812 + j-0.945617675781
            im_multiplicator => "1100001101111011",
            data_re_out => mul_re_out(2004),
            data_im_out => mul_im_out(2004)
        );

 
    UMUL_2005 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2005),
            data_im_in => first_stage_im_out(2005),
            re_multiplicator => "1110010110000111", --- -0.413635253906 + j-0.910461425781
            im_multiplicator => "1100010110111011",
            data_re_out => mul_re_out(2005),
            data_im_out => mul_im_out(2005)
        );

 
    UMUL_2006 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2006),
            data_im_in => first_stage_im_out(2006),
            re_multiplicator => "1110000000011101", --- -0.498229980469 + j-0.867065429688
            im_multiplicator => "1100100010000010",
            data_re_out => mul_re_out(2006),
            data_im_out => mul_im_out(2006)
        );

 
    UMUL_2007 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2007),
            data_im_in => first_stage_im_out(2007),
            re_multiplicator => "1101101011111101", --- -0.578308105469 + j-0.815795898438
            im_multiplicator => "1100101111001010",
            data_re_out => mul_re_out(2007),
            data_im_out => mul_im_out(2007)
        );

 
    UMUL_2008 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2008),
            data_im_in => first_stage_im_out(2008),
            re_multiplicator => "1101011000110010", --- -0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(2008),
            data_im_out => mul_im_out(2008)
        );

 
    UMUL_2009 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2009),
            data_im_in => first_stage_im_out(2009),
            re_multiplicator => "1101000111001001", --- -0.722106933594 + j-0.691772460938
            im_multiplicator => "1101001110111010",
            data_re_out => mul_re_out(2009),
            data_im_out => mul_im_out(2009)
        );

 
    UMUL_2010 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2010),
            data_im_in => first_stage_im_out(2010),
            re_multiplicator => "1100110111001010", --- -0.784545898438 + j-0.620056152344
            im_multiplicator => "1101100001010001",
            data_re_out => mul_re_out(2010),
            data_im_out => mul_im_out(2010)
        );

 
    UMUL_2011 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2011),
            data_im_in => first_stage_im_out(2011),
            re_multiplicator => "1100101000111111", --- -0.839904785156 + j-0.542724609375
            im_multiplicator => "1101110101000100",
            data_re_out => mul_re_out(2011),
            data_im_out => mul_im_out(2011)
        );

 
    UMUL_2012 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2012),
            data_im_in => first_stage_im_out(2012),
            re_multiplicator => "1100011100110001", --- -0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(2012),
            data_im_out => mul_im_out(2012)
        );

 
    UMUL_2013 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2013),
            data_im_in => first_stage_im_out(2013),
            re_multiplicator => "1100010010100110", --- -0.927368164062 + j-0.374145507812
            im_multiplicator => "1110100000001110",
            data_re_out => mul_re_out(2013),
            data_im_out => mul_im_out(2013)
        );

 
    UMUL_2014 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2014),
            data_im_in => first_stage_im_out(2014),
            re_multiplicator => "1100001010100101", --- -0.958679199219 + j-0.284423828125
            im_multiplicator => "1110110111001100",
            data_re_out => mul_re_out(2014),
            data_im_out => mul_im_out(2014)
        );

 
    UMUL_2015 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2015),
            data_im_in => first_stage_im_out(2015),
            re_multiplicator => "1100000100110001", --- -0.981384277344 + j-0.192077636719
            im_multiplicator => "1111001110110101",
            data_re_out => mul_re_out(2015),
            data_im_out => mul_im_out(2015)
        );

 
    UMUL_2016 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2016),
            data_im_in => first_stage_im_out(2016),
            re_multiplicator => "1100000001001111", --- -0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(2016),
            data_im_out => mul_im_out(2016)
        );

 
    UMUL_2017 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2017),
            data_im_in => first_stage_im_out(2017),
            re_multiplicator => "1100000000000000", --- -1.0 + j-0.0030517578125
            im_multiplicator => "1111111111001110",
            data_re_out => mul_re_out(2017),
            data_im_out => mul_im_out(2017)
        );

 
    UMUL_2018 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2018),
            data_im_in => first_stage_im_out(2018),
            re_multiplicator => "1100000001000101", --- -0.995788574219 + j0.0919189453125
            im_multiplicator => "0000010111100010",
            data_re_out => mul_re_out(2018),
            data_im_out => mul_im_out(2018)
        );

 
    UMUL_2019 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2019),
            data_im_in => first_stage_im_out(2019),
            re_multiplicator => "1100000100011110", --- -0.982543945312 + j0.18603515625
            im_multiplicator => "0000101111101000",
            data_re_out => mul_re_out(2019),
            data_im_out => mul_im_out(2019)
        );

 
    UMUL_2020 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2020),
            data_im_in => first_stage_im_out(2020),
            re_multiplicator => "1100001010001000", --- -0.96044921875 + j0.278503417969
            im_multiplicator => "0001000111010011",
            data_re_out => mul_re_out(2020),
            data_im_out => mul_im_out(2020)
        );

 
    UMUL_2021 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2021),
            data_im_in => first_stage_im_out(2021),
            re_multiplicator => "1100010010000001", --- -0.929626464844 + j0.368469238281
            im_multiplicator => "0001011110010101",
            data_re_out => mul_re_out(2021),
            data_im_out => mul_im_out(2021)
        );

 
    UMUL_2022 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2022),
            data_im_in => first_stage_im_out(2022),
            re_multiplicator => "1100011100000011", --- -0.890441894531 + j0.455078125
            im_multiplicator => "0001110100100000",
            data_re_out => mul_re_out(2022),
            data_im_out => mul_im_out(2022)
        );

 
    UMUL_2023 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2023),
            data_im_in => first_stage_im_out(2023),
            re_multiplicator => "1100101000001001", --- -0.843200683594 + j0.53759765625
            im_multiplicator => "0010001001101000",
            data_re_out => mul_re_out(2023),
            data_im_out => mul_im_out(2023)
        );

 
    UMUL_2024 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2024),
            data_im_in => first_stage_im_out(2024),
            re_multiplicator => "1100110110001100", --- -0.788330078125 + j0.615234375
            im_multiplicator => "0010011101100000",
            data_re_out => mul_re_out(2024),
            data_im_out => mul_im_out(2024)
        );

 
    UMUL_2025 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2025),
            data_im_in => first_stage_im_out(2025),
            re_multiplicator => "1101000110000011", --- -0.726379394531 + j0.687316894531
            im_multiplicator => "0010101111111101",
            data_re_out => mul_re_out(2025),
            data_im_out => mul_im_out(2025)
        );

 
    UMUL_2026 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2026),
            data_im_in => first_stage_im_out(2026),
            re_multiplicator => "1101010111100110", --- -0.657836914062 + j0.753173828125
            im_multiplicator => "0011000000110100",
            data_re_out => mul_re_out(2026),
            data_im_out => mul_im_out(2026)
        );

 
    UMUL_2027 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2027),
            data_im_in => first_stage_im_out(2027),
            re_multiplicator => "1101101010101011", --- -0.583312988281 + j0.812255859375
            im_multiplicator => "0011001111111100",
            data_re_out => mul_re_out(2027),
            data_im_out => mul_im_out(2027)
        );

 
    UMUL_2028 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2028),
            data_im_in => first_stage_im_out(2028),
            re_multiplicator => "1101111111000110", --- -0.503540039062 + j0.863952636719
            im_multiplicator => "0011011101001011",
            data_re_out => mul_re_out(2028),
            data_im_out => mul_im_out(2028)
        );

 
    UMUL_2029 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2029),
            data_im_in => first_stage_im_out(2029),
            re_multiplicator => "1110010100101100", --- -0.419189453125 + j0.907897949219
            im_multiplicator => "0011101000011011",
            data_re_out => mul_re_out(2029),
            data_im_out => mul_im_out(2029)
        );

 
    UMUL_2030 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2030),
            data_im_in => first_stage_im_out(2030),
            re_multiplicator => "1110101011001111", --- -0.331115722656 + j0.943603515625
            im_multiplicator => "0011110001100100",
            data_re_out => mul_re_out(2030),
            data_im_out => mul_im_out(2030)
        );

 
    UMUL_2031 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2031),
            data_im_in => first_stage_im_out(2031),
            re_multiplicator => "1111000010100100", --- -0.239990234375 + j0.970764160156
            im_multiplicator => "0011111000100001",
            data_re_out => mul_re_out(2031),
            data_im_out => mul_im_out(2031)
        );

 
    UMUL_2032 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2032),
            data_im_in => first_stage_im_out(2032),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j0.989196777344
            im_multiplicator => "0011111101001111",
            data_re_out => mul_re_out(2032),
            data_im_out => mul_im_out(2032)
        );

 
    UMUL_2033 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2033),
            data_im_in => first_stage_im_out(2033),
            re_multiplicator => "1111110010101010", --- -0.0521240234375 + j0.998657226562
            im_multiplicator => "0011111111101010",
            data_re_out => mul_re_out(2033),
            data_im_out => mul_im_out(2033)
        );

 
    UMUL_2034 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2034),
            data_im_in => first_stage_im_out(2034),
            re_multiplicator => "0000001011000000", --- 0.04296875 + j0.999084472656
            im_multiplicator => "0011111111110001",
            data_re_out => mul_re_out(2034),
            data_im_out => mul_im_out(2034)
        );

 
    UMUL_2035 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2035),
            data_im_in => first_stage_im_out(2035),
            re_multiplicator => "0000100011001111", --- 0.137634277344 + j0.990478515625
            im_multiplicator => "0011111101100100",
            data_re_out => mul_re_out(2035),
            data_im_out => mul_im_out(2035)
        );

 
    UMUL_2036 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2036),
            data_im_in => first_stage_im_out(2036),
            re_multiplicator => "0000111011001010", --- 0.231079101562 + j0.972961425781
            im_multiplicator => "0011111001000101",
            data_re_out => mul_re_out(2036),
            data_im_out => mul_im_out(2036)
        );

 
    UMUL_2037 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2037),
            data_im_in => first_stage_im_out(2037),
            re_multiplicator => "0001010010100010", --- 0.322387695312 + j0.946594238281
            im_multiplicator => "0011110010010101",
            data_re_out => mul_re_out(2037),
            data_im_out => mul_im_out(2037)
        );

 
    UMUL_2038 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2038),
            data_im_in => first_stage_im_out(2038),
            re_multiplicator => "0001101001001011", --- 0.410827636719 + j0.911682128906
            im_multiplicator => "0011101001011001",
            data_re_out => mul_re_out(2038),
            data_im_out => mul_im_out(2038)
        );

 
    UMUL_2039 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2039),
            data_im_in => first_stage_im_out(2039),
            re_multiplicator => "0001111110110111", --- 0.495544433594 + j0.868591308594
            im_multiplicator => "0011011110010111",
            data_re_out => mul_re_out(2039),
            data_im_out => mul_im_out(2039)
        );

 
    UMUL_2040 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2040),
            data_im_in => first_stage_im_out(2040),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j0.817565917969
            im_multiplicator => "0011010001010011",
            data_re_out => mul_re_out(2040),
            data_im_out => mul_im_out(2040)
        );

 
    UMUL_2041 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2041),
            data_im_in => first_stage_im_out(2041),
            re_multiplicator => "0010100110100111", --- 0.650817871094 + j0.759216308594
            im_multiplicator => "0011000010010111",
            data_re_out => mul_re_out(2041),
            data_im_out => mul_im_out(2041)
        );

 
    UMUL_2042 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2042),
            data_im_in => first_stage_im_out(2042),
            re_multiplicator => "0010111000010101", --- 0.720031738281 + j0.693969726562
            im_multiplicator => "0010110001101010",
            data_re_out => mul_re_out(2042),
            data_im_out => mul_im_out(2042)
        );

 
    UMUL_2043 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2043),
            data_im_in => first_stage_im_out(2043),
            re_multiplicator => "0011001000010111", --- 0.782653808594 + j0.622436523438
            im_multiplicator => "0010011111010110",
            data_re_out => mul_re_out(2043),
            data_im_out => mul_im_out(2043)
        );

 
    UMUL_2044 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2044),
            data_im_in => first_stage_im_out(2044),
            re_multiplicator => "0011010110100101", --- 0.838195800781 + j0.545349121094
            im_multiplicator => "0010001011100111",
            data_re_out => mul_re_out(2044),
            data_im_out => mul_im_out(2044)
        );

 
    UMUL_2045 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2045),
            data_im_in => first_stage_im_out(2045),
            re_multiplicator => "0011100010111000", --- 0.88623046875 + j0.463256835938
            im_multiplicator => "0001110110100110",
            data_re_out => mul_re_out(2045),
            data_im_out => mul_im_out(2045)
        );

 
    UMUL_2046 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2046),
            data_im_in => first_stage_im_out(2046),
            re_multiplicator => "0011101101000111", --- 0.926208496094 + j0.377014160156
            im_multiplicator => "0001100000100001",
            data_re_out => mul_re_out(2046),
            data_im_out => mul_im_out(2046)
        );

 
    UMUL_2047 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+5) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(0),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2047),
            data_im_in => first_stage_im_out(2047),
            re_multiplicator => "0011110101001101", --- 0.957824707031 + j0.287353515625
            im_multiplicator => "0001001001100100",
            data_re_out => mul_re_out(2047),
            data_im_out => mul_im_out(2047)
        );

end Behavioral;
