library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity fft_pt512 is
    GENERIC (
        ctrl_start     : INTEGER := 0
    );
    PORT (
        tmp_first_stage_re_out, tmp_first_stage_im_out: OUT STD_LOGIC_VECTOR(511 DOWNTO 0);
        tmp_mul_re_out, tmp_mul_im_out : OUT STD_LOGIC_VECTOR(511 DOWNTO 0);

        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        bypass         : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
        ctrl_delay     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

        data_re_in     : IN STD_LOGIC_VECTOR(511 DOWNTO 0);
        data_im_in     : IN STD_LOGIC_VECTOR(511 DOWNTO 0);

        data_re_out    : OUT STD_LOGIC_VECTOR(511 DOWNTO 0);
        data_im_out    : OUT STD_LOGIC_VECTOR(511 DOWNTO 0)
    );
end fft_pt512;

architecture Behavioral of fft_pt512 is

component fft_pt16 is
    GENERIC (
        ctrl_start     : INTEGER
    );
    PORT (
        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        bypass         : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        ctrl_delay     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

        data_re_in     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_im_in     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

        data_re_out    : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_im_out    : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
end component;

component fft_pt32 is
    GENERIC (
        ctrl_start       : INTEGER
    );
    PORT (
        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        bypass         : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        ctrl_delay     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

        data_re_in     : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        data_im_in     : IN STD_LOGIC_VECTOR(31 DOWNTO 0);

        data_re_out     : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        data_im_out     : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
end component;

component complex_multiplier is
    GENERIC (
        ctrl_start       : INTEGER
    );
    PORT (
        clk              : IN STD_LOGIC;
        rst              : IN STD_LOGIC;
        ce               : IN STD_LOGIC;
        bypass           : IN STD_LOGIC;
        ctrl_delay       : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_in       : IN STD_LOGIC;
        data_im_in       : IN STD_LOGIC;
        re_multiplicator : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        im_multiplicator : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_out      : OUT STD_LOGIC;
        data_im_out      : OUT STD_LOGIC
    );
end component;

component multiplier_mul1 IS
    GENERIC (
        ctrl_start : INTEGER := 0
    );
    PORT (
        clk             : IN STD_LOGIC;
        rst             : IN STD_LOGIC;
        ce              : IN STD_LOGIC;
        bypass          : IN STD_LOGIC;
        ctrl_delay      : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_in      : IN STD_LOGIC;
        data_im_in      : IN STD_LOGIC;
        data_re_out     : OUT STD_LOGIC;
        data_im_out     : OUT STD_LOGIC
    );
END component;

component multiplier_mulminusj IS
    GENERIC (
        ctrl_start : INTEGER := 0
    );
    PORT (
        clk             : IN STD_LOGIC;
        rst             : IN STD_LOGIC;
        ce              : IN STD_LOGIC;
        bypass          : IN STD_LOGIC;
        ctrl_delay      : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_in      : IN STD_LOGIC;
        data_im_in      : IN STD_LOGIC;
        data_re_out     : OUT STD_LOGIC;
        data_im_out     : OUT STD_LOGIC
    );
END component;

COMPONENT Dff_regN_Nout IS
    GENERIC (N : INTEGER);
    PORT (  
        D      : IN STD_LOGIC;
        clk    : IN STD_LOGIC;
        Q      : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        QN     : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0)
    );
END COMPONENT;

--- multiplicator declaration
type ArrOfStdlogic is array (0 to 511) of STD_LOGIC_VECTOR(15 downto 0);
signal re_multiplicator, im_multiplicator : ArrOfStdlogic;

signal first_stage_re_out, first_stage_im_out: STD_LOGIC_VECTOR(511 DOWNTO 0);
signal mul_re_out, mul_im_out : STD_LOGIC_VECTOR(511 DOWNTO 0);

begin
    --- multiplicator definition
    re_multiplicator(33) <= "0011111111111111"; ---  0.999938964844
    im_multiplicator(33) <= "1111111100110111"; --- j-0.0122680664062
    re_multiplicator(34) <= "0011111111111011"; ---  0.999694824219
    im_multiplicator(34) <= "1111111001101110"; --- j-0.0245361328125
    re_multiplicator(35) <= "0011111111110101"; ---  0.999328613281
    im_multiplicator(35) <= "1111110110100101"; --- j-0.0368041992188
    re_multiplicator(36) <= "0011111111101100"; ---  0.998779296875
    im_multiplicator(36) <= "1111110011011100"; --- j-0.049072265625
    re_multiplicator(37) <= "0011111111100001"; ---  0.998107910156
    im_multiplicator(37) <= "1111110000010011"; --- j-0.0613403320312
    re_multiplicator(38) <= "0011111111010100"; ---  0.997314453125
    im_multiplicator(38) <= "1111101101001011"; --- j-0.0735473632812
    re_multiplicator(39) <= "0011111111000100"; ---  0.996337890625
    im_multiplicator(39) <= "1111101010000010"; --- j-0.0858154296875
    re_multiplicator(40) <= "0011111110110001"; ---  0.995178222656
    im_multiplicator(40) <= "1111100110111010"; --- j-0.0980224609375
    re_multiplicator(41) <= "0011111110011100"; ---  0.993896484375
    im_multiplicator(41) <= "1111100011110010"; --- j-0.110229492188
    re_multiplicator(42) <= "0011111110000101"; ---  0.992492675781
    im_multiplicator(42) <= "1111100000101010"; --- j-0.122436523438
    re_multiplicator(43) <= "0011111101101011"; ---  0.990905761719
    im_multiplicator(43) <= "1111011101100011"; --- j-0.134582519531
    re_multiplicator(44) <= "0011111101001111"; ---  0.989196777344
    im_multiplicator(44) <= "1111011010011100"; --- j-0.146728515625
    re_multiplicator(45) <= "0011111100110000"; ---  0.9873046875
    im_multiplicator(45) <= "1111010111010101"; --- j-0.158874511719
    re_multiplicator(46) <= "0011111100001111"; ---  0.985290527344
    im_multiplicator(46) <= "1111010100001111"; --- j-0.170959472656
    re_multiplicator(47) <= "0011111011101011"; ---  0.983093261719
    im_multiplicator(47) <= "1111010001001001"; --- j-0.183044433594
    re_multiplicator(48) <= "0011111011000101"; ---  0.980773925781
    im_multiplicator(48) <= "1111001110000100"; --- j-0.195068359375
    re_multiplicator(49) <= "0011111010011101"; ---  0.978332519531
    im_multiplicator(49) <= "1111001010111111"; --- j-0.207092285156
    re_multiplicator(50) <= "0011111001110010"; ---  0.975708007812
    im_multiplicator(50) <= "1111000111111010"; --- j-0.219116210938
    re_multiplicator(51) <= "0011111001000101"; ---  0.972961425781
    im_multiplicator(51) <= "1111000100110110"; --- j-0.231079101562
    re_multiplicator(52) <= "0011111000010101"; ---  0.970031738281
    im_multiplicator(52) <= "1111000001110011"; --- j-0.242980957031
    re_multiplicator(53) <= "0011110111100011"; ---  0.966979980469
    im_multiplicator(53) <= "1110111110110000"; --- j-0.2548828125
    re_multiplicator(54) <= "0011110110101111"; ---  0.963806152344
    im_multiplicator(54) <= "1110111011101110"; --- j-0.266723632812
    re_multiplicator(55) <= "0011110101111000"; ---  0.96044921875
    im_multiplicator(55) <= "1110111000101101"; --- j-0.278503417969
    re_multiplicator(56) <= "0011110100111111"; ---  0.956970214844
    im_multiplicator(56) <= "1110110101101100"; --- j-0.290283203125
    re_multiplicator(57) <= "0011110100000011"; ---  0.953308105469
    im_multiplicator(57) <= "1110110010101100"; --- j-0.302001953125
    re_multiplicator(58) <= "0011110011000101"; ---  0.949523925781
    im_multiplicator(58) <= "1110101111101101"; --- j-0.313659667969
    re_multiplicator(59) <= "0011110010000101"; ---  0.945617675781
    im_multiplicator(59) <= "1110101100101110"; --- j-0.325317382812
    re_multiplicator(60) <= "0011110001000010"; ---  0.941528320312
    im_multiplicator(60) <= "1110101001110000"; --- j-0.3369140625
    re_multiplicator(61) <= "0011101111111101"; ---  0.937316894531
    im_multiplicator(61) <= "1110100110110100"; --- j-0.348388671875
    re_multiplicator(62) <= "0011101110110110"; ---  0.932983398438
    im_multiplicator(62) <= "1110100011110111"; --- j-0.359924316406
    re_multiplicator(63) <= "0011101101101101"; ---  0.928527832031
    im_multiplicator(63) <= "1110100000111100"; --- j-0.371337890625
    re_multiplicator(65) <= "0011111111111011"; ---  0.999694824219
    im_multiplicator(65) <= "1111111001101110"; --- j-0.0245361328125
    re_multiplicator(66) <= "0011111111101100"; ---  0.998779296875
    im_multiplicator(66) <= "1111110011011100"; --- j-0.049072265625
    re_multiplicator(67) <= "0011111111010100"; ---  0.997314453125
    im_multiplicator(67) <= "1111101101001011"; --- j-0.0735473632812
    re_multiplicator(68) <= "0011111110110001"; ---  0.995178222656
    im_multiplicator(68) <= "1111100110111010"; --- j-0.0980224609375
    re_multiplicator(69) <= "0011111110000101"; ---  0.992492675781
    im_multiplicator(69) <= "1111100000101010"; --- j-0.122436523438
    re_multiplicator(70) <= "0011111101001111"; ---  0.989196777344
    im_multiplicator(70) <= "1111011010011100"; --- j-0.146728515625
    re_multiplicator(71) <= "0011111100001111"; ---  0.985290527344
    im_multiplicator(71) <= "1111010100001111"; --- j-0.170959472656
    re_multiplicator(72) <= "0011111011000101"; ---  0.980773925781
    im_multiplicator(72) <= "1111001110000100"; --- j-0.195068359375
    re_multiplicator(73) <= "0011111001110010"; ---  0.975708007812
    im_multiplicator(73) <= "1111000111111010"; --- j-0.219116210938
    re_multiplicator(74) <= "0011111000010101"; ---  0.970031738281
    im_multiplicator(74) <= "1111000001110011"; --- j-0.242980957031
    re_multiplicator(75) <= "0011110110101111"; ---  0.963806152344
    im_multiplicator(75) <= "1110111011101110"; --- j-0.266723632812
    re_multiplicator(76) <= "0011110100111111"; ---  0.956970214844
    im_multiplicator(76) <= "1110110101101100"; --- j-0.290283203125
    re_multiplicator(77) <= "0011110011000101"; ---  0.949523925781
    im_multiplicator(77) <= "1110101111101101"; --- j-0.313659667969
    re_multiplicator(78) <= "0011110001000010"; ---  0.941528320312
    im_multiplicator(78) <= "1110101001110000"; --- j-0.3369140625
    re_multiplicator(79) <= "0011101110110110"; ---  0.932983398438
    im_multiplicator(79) <= "1110100011110111"; --- j-0.359924316406
    re_multiplicator(80) <= "0011101100100001"; ---  0.923889160156
    im_multiplicator(80) <= "1110011110000010"; --- j-0.382690429688
    re_multiplicator(81) <= "0011101010000010"; ---  0.914184570312
    im_multiplicator(81) <= "1110011000010001"; --- j-0.405212402344
    re_multiplicator(82) <= "0011100111011011"; ---  0.903991699219
    im_multiplicator(82) <= "1110010010100011"; --- j-0.427551269531
    re_multiplicator(83) <= "0011100100101011"; ---  0.893249511719
    im_multiplicator(83) <= "1110001100111010"; --- j-0.449584960938
    re_multiplicator(84) <= "0011100001110001"; ---  0.881896972656
    im_multiplicator(84) <= "1110000111010101"; --- j-0.471374511719
    re_multiplicator(85) <= "0011011110110000"; ---  0.8701171875
    im_multiplicator(85) <= "1110000001110100"; --- j-0.492919921875
    re_multiplicator(86) <= "0011011011100101"; ---  0.857727050781
    im_multiplicator(86) <= "1101111100011001"; --- j-0.514099121094
    re_multiplicator(87) <= "0011011000010010"; ---  0.844848632812
    im_multiplicator(87) <= "1101110111000011"; --- j-0.534973144531
    re_multiplicator(88) <= "0011010100110111"; ---  0.831481933594
    im_multiplicator(88) <= "1101110001110010"; --- j-0.555541992188
    re_multiplicator(89) <= "0011010001010011"; ---  0.817565917969
    im_multiplicator(89) <= "1101101100100110"; --- j-0.575805664062
    re_multiplicator(90) <= "0011001101101000"; ---  0.80322265625
    im_multiplicator(90) <= "1101100111100000"; --- j-0.595703125
    re_multiplicator(91) <= "0011001001110100"; ---  0.788330078125
    im_multiplicator(91) <= "1101100010100000"; --- j-0.615234375
    re_multiplicator(92) <= "0011000101111001"; ---  0.773010253906
    im_multiplicator(92) <= "1101011101100110"; --- j-0.634399414062
    re_multiplicator(93) <= "0011000001110110"; ---  0.757202148438
    im_multiplicator(93) <= "1101011000110010"; --- j-0.653198242188
    re_multiplicator(94) <= "0010111101101100"; ---  0.740966796875
    im_multiplicator(94) <= "1101010100000101"; --- j-0.671569824219
    re_multiplicator(95) <= "0010111001011010"; ---  0.724243164062
    im_multiplicator(95) <= "1101001111011111"; --- j-0.689514160156
    re_multiplicator(97) <= "0011111111110101"; ---  0.999328613281
    im_multiplicator(97) <= "1111110110100101"; --- j-0.0368041992188
    re_multiplicator(98) <= "0011111111010100"; ---  0.997314453125
    im_multiplicator(98) <= "1111101101001011"; --- j-0.0735473632812
    re_multiplicator(99) <= "0011111110011100"; ---  0.993896484375
    im_multiplicator(99) <= "1111100011110010"; --- j-0.110229492188
    re_multiplicator(100) <= "0011111101001111"; ---  0.989196777344
    im_multiplicator(100) <= "1111011010011100"; --- j-0.146728515625
    re_multiplicator(101) <= "0011111011101011"; ---  0.983093261719
    im_multiplicator(101) <= "1111010001001001"; --- j-0.183044433594
    re_multiplicator(102) <= "0011111001110010"; ---  0.975708007812
    im_multiplicator(102) <= "1111000111111010"; --- j-0.219116210938
    re_multiplicator(103) <= "0011110111100011"; ---  0.966979980469
    im_multiplicator(103) <= "1110111110110000"; --- j-0.2548828125
    re_multiplicator(104) <= "0011110100111111"; ---  0.956970214844
    im_multiplicator(104) <= "1110110101101100"; --- j-0.290283203125
    re_multiplicator(105) <= "0011110010000101"; ---  0.945617675781
    im_multiplicator(105) <= "1110101100101110"; --- j-0.325317382812
    re_multiplicator(106) <= "0011101110110110"; ---  0.932983398438
    im_multiplicator(106) <= "1110100011110111"; --- j-0.359924316406
    re_multiplicator(107) <= "0011101011010011"; ---  0.919128417969
    im_multiplicator(107) <= "1110011011001001"; --- j-0.393981933594
    re_multiplicator(108) <= "0011100111011011"; ---  0.903991699219
    im_multiplicator(108) <= "1110010010100011"; --- j-0.427551269531
    re_multiplicator(109) <= "0011100011001111"; ---  0.887634277344
    im_multiplicator(109) <= "1110001010000111"; --- j-0.460510253906
    re_multiplicator(110) <= "0011011110110000"; ---  0.8701171875
    im_multiplicator(110) <= "1110000001110100"; --- j-0.492919921875
    re_multiplicator(111) <= "0011011001111101"; ---  0.851379394531
    im_multiplicator(111) <= "1101111001101101"; --- j-0.524597167969
    re_multiplicator(112) <= "0011010100110111"; ---  0.831481933594
    im_multiplicator(112) <= "1101110001110010"; --- j-0.555541992188
    re_multiplicator(113) <= "0011001111011111"; ---  0.810485839844
    im_multiplicator(113) <= "1101101010000010"; --- j-0.585815429688
    re_multiplicator(114) <= "0011001001110100"; ---  0.788330078125
    im_multiplicator(114) <= "1101100010100000"; --- j-0.615234375
    re_multiplicator(115) <= "0011000011111001"; ---  0.765197753906
    im_multiplicator(115) <= "1101011011001011"; --- j-0.643859863281
    re_multiplicator(116) <= "0010111101101100"; ---  0.740966796875
    im_multiplicator(116) <= "1101010100000101"; --- j-0.671569824219
    re_multiplicator(117) <= "0010110111001111"; ---  0.715759277344
    im_multiplicator(117) <= "1101001101001110"; --- j-0.698364257812
    re_multiplicator(118) <= "0010110000100001"; ---  0.689514160156
    im_multiplicator(118) <= "1101000110100110"; --- j-0.724243164062
    re_multiplicator(119) <= "0010101001100101"; ---  0.662414550781
    im_multiplicator(119) <= "1101000000001110"; --- j-0.749145507812
    re_multiplicator(120) <= "0010100010011010"; ---  0.634399414062
    im_multiplicator(120) <= "1100111010000111"; --- j-0.773010253906
    re_multiplicator(121) <= "0010011011000001"; ---  0.605529785156
    im_multiplicator(121) <= "1100110100010001"; --- j-0.795837402344
    re_multiplicator(122) <= "0010010011011010"; ---  0.575805664062
    im_multiplicator(122) <= "1100101110101101"; --- j-0.817565917969
    re_multiplicator(123) <= "0010001011100111"; ---  0.545349121094
    im_multiplicator(123) <= "1100101001011011"; --- j-0.838195800781
    re_multiplicator(124) <= "0010000011100111"; ---  0.514099121094
    im_multiplicator(124) <= "1100100100011011"; --- j-0.857727050781
    re_multiplicator(125) <= "0001111011011100"; ---  0.482177734375
    im_multiplicator(125) <= "1100011111101110"; --- j-0.876098632812
    re_multiplicator(126) <= "0001110011000110"; ---  0.449584960938
    im_multiplicator(126) <= "1100011011010101"; --- j-0.893249511719
    re_multiplicator(127) <= "0001101010100111"; ---  0.416442871094
    im_multiplicator(127) <= "1100010111010000"; --- j-0.9091796875
    re_multiplicator(129) <= "0011111111101100"; ---  0.998779296875
    im_multiplicator(129) <= "1111110011011100"; --- j-0.049072265625
    re_multiplicator(130) <= "0011111110110001"; ---  0.995178222656
    im_multiplicator(130) <= "1111100110111010"; --- j-0.0980224609375
    re_multiplicator(131) <= "0011111101001111"; ---  0.989196777344
    im_multiplicator(131) <= "1111011010011100"; --- j-0.146728515625
    re_multiplicator(132) <= "0011111011000101"; ---  0.980773925781
    im_multiplicator(132) <= "1111001110000100"; --- j-0.195068359375
    re_multiplicator(133) <= "0011111000010101"; ---  0.970031738281
    im_multiplicator(133) <= "1111000001110011"; --- j-0.242980957031
    re_multiplicator(134) <= "0011110100111111"; ---  0.956970214844
    im_multiplicator(134) <= "1110110101101100"; --- j-0.290283203125
    re_multiplicator(135) <= "0011110001000010"; ---  0.941528320312
    im_multiplicator(135) <= "1110101001110000"; --- j-0.3369140625
    re_multiplicator(136) <= "0011101100100001"; ---  0.923889160156
    im_multiplicator(136) <= "1110011110000010"; --- j-0.382690429688
    re_multiplicator(137) <= "0011100111011011"; ---  0.903991699219
    im_multiplicator(137) <= "1110010010100011"; --- j-0.427551269531
    re_multiplicator(138) <= "0011100001110001"; ---  0.881896972656
    im_multiplicator(138) <= "1110000111010101"; --- j-0.471374511719
    re_multiplicator(139) <= "0011011011100101"; ---  0.857727050781
    im_multiplicator(139) <= "1101111100011001"; --- j-0.514099121094
    re_multiplicator(140) <= "0011010100110111"; ---  0.831481933594
    im_multiplicator(140) <= "1101110001110010"; --- j-0.555541992188
    re_multiplicator(141) <= "0011001101101000"; ---  0.80322265625
    im_multiplicator(141) <= "1101100111100000"; --- j-0.595703125
    re_multiplicator(142) <= "0011000101111001"; ---  0.773010253906
    im_multiplicator(142) <= "1101011101100110"; --- j-0.634399414062
    re_multiplicator(143) <= "0010111101101100"; ---  0.740966796875
    im_multiplicator(143) <= "1101010100000101"; --- j-0.671569824219
    re_multiplicator(144) <= "0010110101000001"; ---  0.707092285156
    im_multiplicator(144) <= "1101001010111111"; --- j-0.707092285156
    re_multiplicator(145) <= "0010101011111011"; ---  0.671569824219
    im_multiplicator(145) <= "1101000010010100"; --- j-0.740966796875
    re_multiplicator(146) <= "0010100010011010"; ---  0.634399414062
    im_multiplicator(146) <= "1100111010000111"; --- j-0.773010253906
    re_multiplicator(147) <= "0010011000100000"; ---  0.595703125
    im_multiplicator(147) <= "1100110010011000"; --- j-0.80322265625
    re_multiplicator(148) <= "0010001110001110"; ---  0.555541992188
    im_multiplicator(148) <= "1100101011001001"; --- j-0.831481933594
    re_multiplicator(149) <= "0010000011100111"; ---  0.514099121094
    im_multiplicator(149) <= "1100100100011011"; --- j-0.857727050781
    re_multiplicator(150) <= "0001111000101011"; ---  0.471374511719
    im_multiplicator(150) <= "1100011110001111"; --- j-0.881896972656
    re_multiplicator(151) <= "0001101101011101"; ---  0.427551269531
    im_multiplicator(151) <= "1100011000100101"; --- j-0.903991699219
    re_multiplicator(152) <= "0001100001111110"; ---  0.382690429688
    im_multiplicator(152) <= "1100010011011111"; --- j-0.923889160156
    re_multiplicator(153) <= "0001010110010000"; ---  0.3369140625
    im_multiplicator(153) <= "1100001110111110"; --- j-0.941528320312
    re_multiplicator(154) <= "0001001010010100"; ---  0.290283203125
    im_multiplicator(154) <= "1100001011000001"; --- j-0.956970214844
    re_multiplicator(155) <= "0000111110001101"; ---  0.242980957031
    im_multiplicator(155) <= "1100000111101011"; --- j-0.970031738281
    re_multiplicator(156) <= "0000110001111100"; ---  0.195068359375
    im_multiplicator(156) <= "1100000100111011"; --- j-0.980773925781
    re_multiplicator(157) <= "0000100101100100"; ---  0.146728515625
    im_multiplicator(157) <= "1100000010110001"; --- j-0.989196777344
    re_multiplicator(158) <= "0000011001000110"; ---  0.0980224609375
    im_multiplicator(158) <= "1100000001001111"; --- j-0.995178222656
    re_multiplicator(159) <= "0000001100100100"; ---  0.049072265625
    im_multiplicator(159) <= "1100000000010100"; --- j-0.998779296875
    re_multiplicator(161) <= "0011111111100001"; ---  0.998107910156
    im_multiplicator(161) <= "1111110000010011"; --- j-0.0613403320312
    re_multiplicator(162) <= "0011111110000101"; ---  0.992492675781
    im_multiplicator(162) <= "1111100000101010"; --- j-0.122436523438
    re_multiplicator(163) <= "0011111011101011"; ---  0.983093261719
    im_multiplicator(163) <= "1111010001001001"; --- j-0.183044433594
    re_multiplicator(164) <= "0011111000010101"; ---  0.970031738281
    im_multiplicator(164) <= "1111000001110011"; --- j-0.242980957031
    re_multiplicator(165) <= "0011110100000011"; ---  0.953308105469
    im_multiplicator(165) <= "1110110010101100"; --- j-0.302001953125
    re_multiplicator(166) <= "0011101110110110"; ---  0.932983398438
    im_multiplicator(166) <= "1110100011110111"; --- j-0.359924316406
    re_multiplicator(167) <= "0011101000110000"; ---  0.9091796875
    im_multiplicator(167) <= "1110010101011001"; --- j-0.416442871094
    re_multiplicator(168) <= "0011100001110001"; ---  0.881896972656
    im_multiplicator(168) <= "1110000111010101"; --- j-0.471374511719
    re_multiplicator(169) <= "0011011001111101"; ---  0.851379394531
    im_multiplicator(169) <= "1101111001101101"; --- j-0.524597167969
    re_multiplicator(170) <= "0011010001010011"; ---  0.817565917969
    im_multiplicator(170) <= "1101101100100110"; --- j-0.575805664062
    re_multiplicator(171) <= "0011000111111000"; ---  0.78076171875
    im_multiplicator(171) <= "1101100000000010"; --- j-0.624877929688
    re_multiplicator(172) <= "0010111101101100"; ---  0.740966796875
    im_multiplicator(172) <= "1101010100000101"; --- j-0.671569824219
    re_multiplicator(173) <= "0010110010110010"; ---  0.698364257812
    im_multiplicator(173) <= "1101001000110001"; --- j-0.715759277344
    re_multiplicator(174) <= "0010100111001110"; ---  0.653198242188
    im_multiplicator(174) <= "1100111110001010"; --- j-0.757202148438
    re_multiplicator(175) <= "0010011011000001"; ---  0.605529785156
    im_multiplicator(175) <= "1100110100010001"; --- j-0.795837402344
    re_multiplicator(176) <= "0010001110001110"; ---  0.555541992188
    im_multiplicator(176) <= "1100101011001001"; --- j-0.831481933594
    re_multiplicator(177) <= "0010000000111010"; ---  0.503540039062
    im_multiplicator(177) <= "1100100010110101"; --- j-0.863952636719
    re_multiplicator(178) <= "0001110011000110"; ---  0.449584960938
    im_multiplicator(178) <= "1100011011010101"; --- j-0.893249511719
    re_multiplicator(179) <= "0001100100110111"; ---  0.393981933594
    im_multiplicator(179) <= "1100010100101101"; --- j-0.919128417969
    re_multiplicator(180) <= "0001010110010000"; ---  0.3369140625
    im_multiplicator(180) <= "1100001110111110"; --- j-0.941528320312
    re_multiplicator(181) <= "0001000111010011"; ---  0.278503417969
    im_multiplicator(181) <= "1100001010001000"; --- j-0.96044921875
    re_multiplicator(182) <= "0000111000000110"; ---  0.219116210938
    im_multiplicator(182) <= "1100000110001110"; --- j-0.975708007812
    re_multiplicator(183) <= "0000101000101011"; ---  0.158874511719
    im_multiplicator(183) <= "1100000011010000"; --- j-0.9873046875
    re_multiplicator(184) <= "0000011001000110"; ---  0.0980224609375
    im_multiplicator(184) <= "1100000001001111"; --- j-0.995178222656
    re_multiplicator(185) <= "0000001001011011"; ---  0.0368041992188
    im_multiplicator(185) <= "1100000000001011"; --- j-0.999328613281
    re_multiplicator(186) <= "1111111001101110"; ---  -0.0245361328125
    im_multiplicator(186) <= "1100000000000101"; --- j-0.999694824219
    re_multiplicator(187) <= "1111101010000010"; ---  -0.0858154296875
    im_multiplicator(187) <= "1100000000111100"; --- j-0.996337890625
    re_multiplicator(188) <= "1111011010011100"; ---  -0.146728515625
    im_multiplicator(188) <= "1100000010110001"; --- j-0.989196777344
    re_multiplicator(189) <= "1111001010111111"; ---  -0.207092285156
    im_multiplicator(189) <= "1100000101100011"; --- j-0.978332519531
    re_multiplicator(190) <= "1110111011101110"; ---  -0.266723632812
    im_multiplicator(190) <= "1100001001010001"; --- j-0.963806152344
    re_multiplicator(191) <= "1110101100101110"; ---  -0.325317382812
    im_multiplicator(191) <= "1100001101111011"; --- j-0.945617675781
    re_multiplicator(193) <= "0011111111010100"; ---  0.997314453125
    im_multiplicator(193) <= "1111101101001011"; --- j-0.0735473632812
    re_multiplicator(194) <= "0011111101001111"; ---  0.989196777344
    im_multiplicator(194) <= "1111011010011100"; --- j-0.146728515625
    re_multiplicator(195) <= "0011111001110010"; ---  0.975708007812
    im_multiplicator(195) <= "1111000111111010"; --- j-0.219116210938
    re_multiplicator(196) <= "0011110100111111"; ---  0.956970214844
    im_multiplicator(196) <= "1110110101101100"; --- j-0.290283203125
    re_multiplicator(197) <= "0011101110110110"; ---  0.932983398438
    im_multiplicator(197) <= "1110100011110111"; --- j-0.359924316406
    re_multiplicator(198) <= "0011100111011011"; ---  0.903991699219
    im_multiplicator(198) <= "1110010010100011"; --- j-0.427551269531
    re_multiplicator(199) <= "0011011110110000"; ---  0.8701171875
    im_multiplicator(199) <= "1110000001110100"; --- j-0.492919921875
    re_multiplicator(200) <= "0011010100110111"; ---  0.831481933594
    im_multiplicator(200) <= "1101110001110010"; --- j-0.555541992188
    re_multiplicator(201) <= "0011001001110100"; ---  0.788330078125
    im_multiplicator(201) <= "1101100010100000"; --- j-0.615234375
    re_multiplicator(202) <= "0010111101101100"; ---  0.740966796875
    im_multiplicator(202) <= "1101010100000101"; --- j-0.671569824219
    re_multiplicator(203) <= "0010110000100001"; ---  0.689514160156
    im_multiplicator(203) <= "1101000110100110"; --- j-0.724243164062
    re_multiplicator(204) <= "0010100010011010"; ---  0.634399414062
    im_multiplicator(204) <= "1100111010000111"; --- j-0.773010253906
    re_multiplicator(205) <= "0010010011011010"; ---  0.575805664062
    im_multiplicator(205) <= "1100101110101101"; --- j-0.817565917969
    re_multiplicator(206) <= "0010000011100111"; ---  0.514099121094
    im_multiplicator(206) <= "1100100100011011"; --- j-0.857727050781
    re_multiplicator(207) <= "0001110011000110"; ---  0.449584960938
    im_multiplicator(207) <= "1100011011010101"; --- j-0.893249511719
    re_multiplicator(208) <= "0001100001111110"; ---  0.382690429688
    im_multiplicator(208) <= "1100010011011111"; --- j-0.923889160156
    re_multiplicator(209) <= "0001010000010011"; ---  0.313659667969
    im_multiplicator(209) <= "1100001100111011"; --- j-0.949523925781
    re_multiplicator(210) <= "0000111110001101"; ---  0.242980957031
    im_multiplicator(210) <= "1100000111101011"; --- j-0.970031738281
    re_multiplicator(211) <= "0000101011110001"; ---  0.170959472656
    im_multiplicator(211) <= "1100000011110001"; --- j-0.985290527344
    re_multiplicator(212) <= "0000011001000110"; ---  0.0980224609375
    im_multiplicator(212) <= "1100000001001111"; --- j-0.995178222656
    re_multiplicator(213) <= "0000000110010010"; ---  0.0245361328125
    im_multiplicator(213) <= "1100000000000101"; --- j-0.999694824219
    re_multiplicator(214) <= "1111110011011100"; ---  -0.049072265625
    im_multiplicator(214) <= "1100000000010100"; --- j-0.998779296875
    re_multiplicator(215) <= "1111100000101010"; ---  -0.122436523438
    im_multiplicator(215) <= "1100000001111011"; --- j-0.992492675781
    re_multiplicator(216) <= "1111001110000100"; ---  -0.195068359375
    im_multiplicator(216) <= "1100000100111011"; --- j-0.980773925781
    re_multiplicator(217) <= "1110111011101110"; ---  -0.266723632812
    im_multiplicator(217) <= "1100001001010001"; --- j-0.963806152344
    re_multiplicator(218) <= "1110101001110000"; ---  -0.3369140625
    im_multiplicator(218) <= "1100001110111110"; --- j-0.941528320312
    re_multiplicator(219) <= "1110011000010001"; ---  -0.405212402344
    im_multiplicator(219) <= "1100010101111110"; --- j-0.914184570312
    re_multiplicator(220) <= "1110000111010101"; ---  -0.471374511719
    im_multiplicator(220) <= "1100011110001111"; --- j-0.881896972656
    re_multiplicator(221) <= "1101110111000011"; ---  -0.534973144531
    im_multiplicator(221) <= "1100100111101110"; --- j-0.844848632812
    re_multiplicator(222) <= "1101100111100000"; ---  -0.595703125
    im_multiplicator(222) <= "1100110010011000"; --- j-0.80322265625
    re_multiplicator(223) <= "1101011000110010"; ---  -0.653198242188
    im_multiplicator(223) <= "1100111110001010"; --- j-0.757202148438
    re_multiplicator(225) <= "0011111111000100"; ---  0.996337890625
    im_multiplicator(225) <= "1111101010000010"; --- j-0.0858154296875
    re_multiplicator(226) <= "0011111100001111"; ---  0.985290527344
    im_multiplicator(226) <= "1111010100001111"; --- j-0.170959472656
    re_multiplicator(227) <= "0011110111100011"; ---  0.966979980469
    im_multiplicator(227) <= "1110111110110000"; --- j-0.2548828125
    re_multiplicator(228) <= "0011110001000010"; ---  0.941528320312
    im_multiplicator(228) <= "1110101001110000"; --- j-0.3369140625
    re_multiplicator(229) <= "0011101000110000"; ---  0.9091796875
    im_multiplicator(229) <= "1110010101011001"; --- j-0.416442871094
    re_multiplicator(230) <= "0011011110110000"; ---  0.8701171875
    im_multiplicator(230) <= "1110000001110100"; --- j-0.492919921875
    re_multiplicator(231) <= "0011010011000110"; ---  0.824584960938
    im_multiplicator(231) <= "1101101111001011"; --- j-0.565734863281
    re_multiplicator(232) <= "0011000101111001"; ---  0.773010253906
    im_multiplicator(232) <= "1101011101100110"; --- j-0.634399414062
    re_multiplicator(233) <= "0010110111001111"; ---  0.715759277344
    im_multiplicator(233) <= "1101001101001110"; --- j-0.698364257812
    re_multiplicator(234) <= "0010100111001110"; ---  0.653198242188
    im_multiplicator(234) <= "1100111110001010"; --- j-0.757202148438
    re_multiplicator(235) <= "0010010101111110"; ---  0.585815429688
    im_multiplicator(235) <= "1100110000100001"; --- j-0.810485839844
    re_multiplicator(236) <= "0010000011100111"; ---  0.514099121094
    im_multiplicator(236) <= "1100100100011011"; --- j-0.857727050781
    re_multiplicator(237) <= "0001110000010010"; ---  0.438598632812
    im_multiplicator(237) <= "1100011001111100"; --- j-0.898681640625
    re_multiplicator(238) <= "0001011100001001"; ---  0.359924316406
    im_multiplicator(238) <= "1100010001001010"; --- j-0.932983398438
    re_multiplicator(239) <= "0001000111010011"; ---  0.278503417969
    im_multiplicator(239) <= "1100001010001000"; --- j-0.96044921875
    re_multiplicator(240) <= "0000110001111100"; ---  0.195068359375
    im_multiplicator(240) <= "1100000100111011"; --- j-0.980773925781
    re_multiplicator(241) <= "0000011100001110"; ---  0.110229492188
    im_multiplicator(241) <= "1100000001100100"; --- j-0.993896484375
    re_multiplicator(242) <= "0000000110010010"; ---  0.0245361328125
    im_multiplicator(242) <= "1100000000000101"; --- j-0.999694824219
    re_multiplicator(243) <= "1111110000010011"; ---  -0.0613403320312
    im_multiplicator(243) <= "1100000000011111"; --- j-0.998107910156
    re_multiplicator(244) <= "1111011010011100"; ---  -0.146728515625
    im_multiplicator(244) <= "1100000010110001"; --- j-0.989196777344
    re_multiplicator(245) <= "1111000100110110"; ---  -0.231079101562
    im_multiplicator(245) <= "1100000110111011"; --- j-0.972961425781
    re_multiplicator(246) <= "1110101111101101"; ---  -0.313659667969
    im_multiplicator(246) <= "1100001100111011"; --- j-0.949523925781
    re_multiplicator(247) <= "1110011011001001"; ---  -0.393981933594
    im_multiplicator(247) <= "1100010100101101"; --- j-0.919128417969
    re_multiplicator(248) <= "1110000111010101"; ---  -0.471374511719
    im_multiplicator(248) <= "1100011110001111"; --- j-0.881896972656
    re_multiplicator(249) <= "1101110100011001"; ---  -0.545349121094
    im_multiplicator(249) <= "1100101001011011"; --- j-0.838195800781
    re_multiplicator(250) <= "1101100010100000"; ---  -0.615234375
    im_multiplicator(250) <= "1100110110001100"; --- j-0.788330078125
    re_multiplicator(251) <= "1101010001110001"; ---  -0.680603027344
    im_multiplicator(251) <= "1101000100011100"; --- j-0.732666015625
    re_multiplicator(252) <= "1101000010010100"; ---  -0.740966796875
    im_multiplicator(252) <= "1101010100000101"; --- j-0.671569824219
    re_multiplicator(253) <= "1100110100010001"; ---  -0.795837402344
    im_multiplicator(253) <= "1101100100111111"; --- j-0.605529785156
    re_multiplicator(254) <= "1100100111101110"; ---  -0.844848632812
    im_multiplicator(254) <= "1101110111000011"; --- j-0.534973144531
    re_multiplicator(255) <= "1100011100110001"; ---  -0.887634277344
    im_multiplicator(255) <= "1110001010000111"; --- j-0.460510253906
    re_multiplicator(257) <= "0011111110110001"; ---  0.995178222656
    im_multiplicator(257) <= "1111100110111010"; --- j-0.0980224609375
    re_multiplicator(258) <= "0011111011000101"; ---  0.980773925781
    im_multiplicator(258) <= "1111001110000100"; --- j-0.195068359375
    re_multiplicator(259) <= "0011110100111111"; ---  0.956970214844
    im_multiplicator(259) <= "1110110101101100"; --- j-0.290283203125
    re_multiplicator(260) <= "0011101100100001"; ---  0.923889160156
    im_multiplicator(260) <= "1110011110000010"; --- j-0.382690429688
    re_multiplicator(261) <= "0011100001110001"; ---  0.881896972656
    im_multiplicator(261) <= "1110000111010101"; --- j-0.471374511719
    re_multiplicator(262) <= "0011010100110111"; ---  0.831481933594
    im_multiplicator(262) <= "1101110001110010"; --- j-0.555541992188
    re_multiplicator(263) <= "0011000101111001"; ---  0.773010253906
    im_multiplicator(263) <= "1101011101100110"; --- j-0.634399414062
    re_multiplicator(264) <= "0010110101000001"; ---  0.707092285156
    im_multiplicator(264) <= "1101001010111111"; --- j-0.707092285156
    re_multiplicator(265) <= "0010100010011010"; ---  0.634399414062
    im_multiplicator(265) <= "1100111010000111"; --- j-0.773010253906
    re_multiplicator(266) <= "0010001110001110"; ---  0.555541992188
    im_multiplicator(266) <= "1100101011001001"; --- j-0.831481933594
    re_multiplicator(267) <= "0001111000101011"; ---  0.471374511719
    im_multiplicator(267) <= "1100011110001111"; --- j-0.881896972656
    re_multiplicator(268) <= "0001100001111110"; ---  0.382690429688
    im_multiplicator(268) <= "1100010011011111"; --- j-0.923889160156
    re_multiplicator(269) <= "0001001010010100"; ---  0.290283203125
    im_multiplicator(269) <= "1100001011000001"; --- j-0.956970214844
    re_multiplicator(270) <= "0000110001111100"; ---  0.195068359375
    im_multiplicator(270) <= "1100000100111011"; --- j-0.980773925781
    re_multiplicator(271) <= "0000011001000110"; ---  0.0980224609375
    im_multiplicator(271) <= "1100000001001111"; --- j-0.995178222656
    re_multiplicator(273) <= "1111100110111010"; ---  -0.0980224609375
    im_multiplicator(273) <= "1100000001001111"; --- j-0.995178222656
    re_multiplicator(274) <= "1111001110000100"; ---  -0.195068359375
    im_multiplicator(274) <= "1100000100111011"; --- j-0.980773925781
    re_multiplicator(275) <= "1110110101101100"; ---  -0.290283203125
    im_multiplicator(275) <= "1100001011000001"; --- j-0.956970214844
    re_multiplicator(276) <= "1110011110000010"; ---  -0.382690429688
    im_multiplicator(276) <= "1100010011011111"; --- j-0.923889160156
    re_multiplicator(277) <= "1110000111010101"; ---  -0.471374511719
    im_multiplicator(277) <= "1100011110001111"; --- j-0.881896972656
    re_multiplicator(278) <= "1101110001110010"; ---  -0.555541992188
    im_multiplicator(278) <= "1100101011001001"; --- j-0.831481933594
    re_multiplicator(279) <= "1101011101100110"; ---  -0.634399414062
    im_multiplicator(279) <= "1100111010000111"; --- j-0.773010253906
    re_multiplicator(280) <= "1101001010111111"; ---  -0.707092285156
    im_multiplicator(280) <= "1101001010111111"; --- j-0.707092285156
    re_multiplicator(281) <= "1100111010000111"; ---  -0.773010253906
    im_multiplicator(281) <= "1101011101100110"; --- j-0.634399414062
    re_multiplicator(282) <= "1100101011001001"; ---  -0.831481933594
    im_multiplicator(282) <= "1101110001110010"; --- j-0.555541992188
    re_multiplicator(283) <= "1100011110001111"; ---  -0.881896972656
    im_multiplicator(283) <= "1110000111010101"; --- j-0.471374511719
    re_multiplicator(284) <= "1100010011011111"; ---  -0.923889160156
    im_multiplicator(284) <= "1110011110000010"; --- j-0.382690429688
    re_multiplicator(285) <= "1100001011000001"; ---  -0.956970214844
    im_multiplicator(285) <= "1110110101101100"; --- j-0.290283203125
    re_multiplicator(286) <= "1100000100111011"; ---  -0.980773925781
    im_multiplicator(286) <= "1111001110000100"; --- j-0.195068359375
    re_multiplicator(287) <= "1100000001001111"; ---  -0.995178222656
    im_multiplicator(287) <= "1111100110111010"; --- j-0.0980224609375
    re_multiplicator(289) <= "0011111110011100"; ---  0.993896484375
    im_multiplicator(289) <= "1111100011110010"; --- j-0.110229492188
    re_multiplicator(290) <= "0011111001110010"; ---  0.975708007812
    im_multiplicator(290) <= "1111000111111010"; --- j-0.219116210938
    re_multiplicator(291) <= "0011110010000101"; ---  0.945617675781
    im_multiplicator(291) <= "1110101100101110"; --- j-0.325317382812
    re_multiplicator(292) <= "0011100111011011"; ---  0.903991699219
    im_multiplicator(292) <= "1110010010100011"; --- j-0.427551269531
    re_multiplicator(293) <= "0011011001111101"; ---  0.851379394531
    im_multiplicator(293) <= "1101111001101101"; --- j-0.524597167969
    re_multiplicator(294) <= "0011001001110100"; ---  0.788330078125
    im_multiplicator(294) <= "1101100010100000"; --- j-0.615234375
    re_multiplicator(295) <= "0010110111001111"; ---  0.715759277344
    im_multiplicator(295) <= "1101001101001110"; --- j-0.698364257812
    re_multiplicator(296) <= "0010100010011010"; ---  0.634399414062
    im_multiplicator(296) <= "1100111010000111"; --- j-0.773010253906
    re_multiplicator(297) <= "0010001011100111"; ---  0.545349121094
    im_multiplicator(297) <= "1100101001011011"; --- j-0.838195800781
    re_multiplicator(298) <= "0001110011000110"; ---  0.449584960938
    im_multiplicator(298) <= "1100011011010101"; --- j-0.893249511719
    re_multiplicator(299) <= "0001011001001100"; ---  0.348388671875
    im_multiplicator(299) <= "1100010000000011"; --- j-0.937316894531
    re_multiplicator(300) <= "0000111110001101"; ---  0.242980957031
    im_multiplicator(300) <= "1100000111101011"; --- j-0.970031738281
    re_multiplicator(301) <= "0000100010011101"; ---  0.134582519531
    im_multiplicator(301) <= "1100000010010101"; --- j-0.990905761719
    re_multiplicator(302) <= "0000000110010010"; ---  0.0245361328125
    im_multiplicator(302) <= "1100000000000101"; --- j-0.999694824219
    re_multiplicator(303) <= "1111101010000010"; ---  -0.0858154296875
    im_multiplicator(303) <= "1100000000111100"; --- j-0.996337890625
    re_multiplicator(304) <= "1111001110000100"; ---  -0.195068359375
    im_multiplicator(304) <= "1100000100111011"; --- j-0.980773925781
    re_multiplicator(305) <= "1110110010101100"; ---  -0.302001953125
    im_multiplicator(305) <= "1100001011111101"; --- j-0.953308105469
    re_multiplicator(306) <= "1110011000010001"; ---  -0.405212402344
    im_multiplicator(306) <= "1100010101111110"; --- j-0.914184570312
    re_multiplicator(307) <= "1101111111000110"; ---  -0.503540039062
    im_multiplicator(307) <= "1100100010110101"; --- j-0.863952636719
    re_multiplicator(308) <= "1101100111100000"; ---  -0.595703125
    im_multiplicator(308) <= "1100110010011000"; --- j-0.80322265625
    re_multiplicator(309) <= "1101010001110001"; ---  -0.680603027344
    im_multiplicator(309) <= "1101000100011100"; --- j-0.732666015625
    re_multiplicator(310) <= "1100111110001010"; ---  -0.757202148438
    im_multiplicator(310) <= "1101011000110010"; --- j-0.653198242188
    re_multiplicator(311) <= "1100101100111010"; ---  -0.824584960938
    im_multiplicator(311) <= "1101101111001011"; --- j-0.565734863281
    re_multiplicator(312) <= "1100011110001111"; ---  -0.881896972656
    im_multiplicator(312) <= "1110000111010101"; --- j-0.471374511719
    re_multiplicator(313) <= "1100010010010011"; ---  -0.928527832031
    im_multiplicator(313) <= "1110100000111100"; --- j-0.371337890625
    re_multiplicator(314) <= "1100001001010001"; ---  -0.963806152344
    im_multiplicator(314) <= "1110111011101110"; --- j-0.266723632812
    re_multiplicator(315) <= "1100000011010000"; ---  -0.9873046875
    im_multiplicator(315) <= "1111010111010101"; --- j-0.158874511719
    re_multiplicator(316) <= "1100000000010100"; ---  -0.998779296875
    im_multiplicator(316) <= "1111110011011100"; --- j-0.049072265625
    re_multiplicator(317) <= "1100000000011111"; ---  -0.998107910156
    im_multiplicator(317) <= "0000001111101101"; --- j0.0613403320312
    re_multiplicator(318) <= "1100000011110001"; ---  -0.985290527344
    im_multiplicator(318) <= "0000101011110001"; --- j0.170959472656
    re_multiplicator(319) <= "1100001010001000"; ---  -0.96044921875
    im_multiplicator(319) <= "0001000111010011"; --- j0.278503417969
    re_multiplicator(321) <= "0011111110000101"; ---  0.992492675781
    im_multiplicator(321) <= "1111100000101010"; --- j-0.122436523438
    re_multiplicator(322) <= "0011111000010101"; ---  0.970031738281
    im_multiplicator(322) <= "1111000001110011"; --- j-0.242980957031
    re_multiplicator(323) <= "0011101110110110"; ---  0.932983398438
    im_multiplicator(323) <= "1110100011110111"; --- j-0.359924316406
    re_multiplicator(324) <= "0011100001110001"; ---  0.881896972656
    im_multiplicator(324) <= "1110000111010101"; --- j-0.471374511719
    re_multiplicator(325) <= "0011010001010011"; ---  0.817565917969
    im_multiplicator(325) <= "1101101100100110"; --- j-0.575805664062
    re_multiplicator(326) <= "0010111101101100"; ---  0.740966796875
    im_multiplicator(326) <= "1101010100000101"; --- j-0.671569824219
    re_multiplicator(327) <= "0010100111001110"; ---  0.653198242188
    im_multiplicator(327) <= "1100111110001010"; --- j-0.757202148438
    re_multiplicator(328) <= "0010001110001110"; ---  0.555541992188
    im_multiplicator(328) <= "1100101011001001"; --- j-0.831481933594
    re_multiplicator(329) <= "0001110011000110"; ---  0.449584960938
    im_multiplicator(329) <= "1100011011010101"; --- j-0.893249511719
    re_multiplicator(330) <= "0001010110010000"; ---  0.3369140625
    im_multiplicator(330) <= "1100001110111110"; --- j-0.941528320312
    re_multiplicator(331) <= "0000111000000110"; ---  0.219116210938
    im_multiplicator(331) <= "1100000110001110"; --- j-0.975708007812
    re_multiplicator(332) <= "0000011001000110"; ---  0.0980224609375
    im_multiplicator(332) <= "1100000001001111"; --- j-0.995178222656
    re_multiplicator(333) <= "1111111001101110"; ---  -0.0245361328125
    im_multiplicator(333) <= "1100000000000101"; --- j-0.999694824219
    re_multiplicator(334) <= "1111011010011100"; ---  -0.146728515625
    im_multiplicator(334) <= "1100000010110001"; --- j-0.989196777344
    re_multiplicator(335) <= "1110111011101110"; ---  -0.266723632812
    im_multiplicator(335) <= "1100001001010001"; --- j-0.963806152344
    re_multiplicator(336) <= "1110011110000010"; ---  -0.382690429688
    im_multiplicator(336) <= "1100010011011111"; --- j-0.923889160156
    re_multiplicator(337) <= "1110000001110100"; ---  -0.492919921875
    im_multiplicator(337) <= "1100100001010000"; --- j-0.8701171875
    re_multiplicator(338) <= "1101100111100000"; ---  -0.595703125
    im_multiplicator(338) <= "1100110010011000"; --- j-0.80322265625
    re_multiplicator(339) <= "1101001111011111"; ---  -0.689514160156
    im_multiplicator(339) <= "1101000110100110"; --- j-0.724243164062
    re_multiplicator(340) <= "1100111010000111"; ---  -0.773010253906
    im_multiplicator(340) <= "1101011101100110"; --- j-0.634399414062
    re_multiplicator(341) <= "1100100111101110"; ---  -0.844848632812
    im_multiplicator(341) <= "1101110111000011"; --- j-0.534973144531
    re_multiplicator(342) <= "1100011000100101"; ---  -0.903991699219
    im_multiplicator(342) <= "1110010010100011"; --- j-0.427551269531
    re_multiplicator(343) <= "1100001100111011"; ---  -0.949523925781
    im_multiplicator(343) <= "1110101111101101"; --- j-0.313659667969
    re_multiplicator(344) <= "1100000100111011"; ---  -0.980773925781
    im_multiplicator(344) <= "1111001110000100"; --- j-0.195068359375
    re_multiplicator(345) <= "1100000000101100"; ---  -0.997314453125
    im_multiplicator(345) <= "1111101101001011"; --- j-0.0735473632812
    re_multiplicator(346) <= "1100000000010100"; ---  -0.998779296875
    im_multiplicator(346) <= "0000001100100100"; --- j0.049072265625
    re_multiplicator(347) <= "1100000011110001"; ---  -0.985290527344
    im_multiplicator(347) <= "0000101011110001"; --- j0.170959472656
    re_multiplicator(348) <= "1100001011000001"; ---  -0.956970214844
    im_multiplicator(348) <= "0001001010010100"; --- j0.290283203125
    re_multiplicator(349) <= "1100010101111110"; ---  -0.914184570312
    im_multiplicator(349) <= "0001100111101111"; --- j0.405212402344
    re_multiplicator(350) <= "1100100100011011"; ---  -0.857727050781
    im_multiplicator(350) <= "0010000011100111"; --- j0.514099121094
    re_multiplicator(351) <= "1100110110001100"; ---  -0.788330078125
    im_multiplicator(351) <= "0010011101100000"; --- j0.615234375
    re_multiplicator(353) <= "0011111101101011"; ---  0.990905761719
    im_multiplicator(353) <= "1111011101100011"; --- j-0.134582519531
    re_multiplicator(354) <= "0011110110101111"; ---  0.963806152344
    im_multiplicator(354) <= "1110111011101110"; --- j-0.266723632812
    re_multiplicator(355) <= "0011101011010011"; ---  0.919128417969
    im_multiplicator(355) <= "1110011011001001"; --- j-0.393981933594
    re_multiplicator(356) <= "0011011011100101"; ---  0.857727050781
    im_multiplicator(356) <= "1101111100011001"; --- j-0.514099121094
    re_multiplicator(357) <= "0011000111111000"; ---  0.78076171875
    im_multiplicator(357) <= "1101100000000010"; --- j-0.624877929688
    re_multiplicator(358) <= "0010110000100001"; ---  0.689514160156
    im_multiplicator(358) <= "1101000110100110"; --- j-0.724243164062
    re_multiplicator(359) <= "0010010101111110"; ---  0.585815429688
    im_multiplicator(359) <= "1100110000100001"; --- j-0.810485839844
    re_multiplicator(360) <= "0001111000101011"; ---  0.471374511719
    im_multiplicator(360) <= "1100011110001111"; --- j-0.881896972656
    re_multiplicator(361) <= "0001011001001100"; ---  0.348388671875
    im_multiplicator(361) <= "1100010000000011"; --- j-0.937316894531
    re_multiplicator(362) <= "0000111000000110"; ---  0.219116210938
    im_multiplicator(362) <= "1100000110001110"; --- j-0.975708007812
    re_multiplicator(363) <= "0000010101111110"; ---  0.0858154296875
    im_multiplicator(363) <= "1100000000111100"; --- j-0.996337890625
    re_multiplicator(364) <= "1111110011011100"; ---  -0.049072265625
    im_multiplicator(364) <= "1100000000010100"; --- j-0.998779296875
    re_multiplicator(365) <= "1111010001001001"; ---  -0.183044433594
    im_multiplicator(365) <= "1100000100010101"; --- j-0.983093261719
    re_multiplicator(366) <= "1110101111101101"; ---  -0.313659667969
    im_multiplicator(366) <= "1100001100111011"; --- j-0.949523925781
    re_multiplicator(367) <= "1110001111101110"; ---  -0.438598632812
    im_multiplicator(367) <= "1100011001111100"; --- j-0.898681640625
    re_multiplicator(368) <= "1101110001110010"; ---  -0.555541992188
    im_multiplicator(368) <= "1100101011001001"; --- j-0.831481933594
    re_multiplicator(369) <= "1101010110011011"; ---  -0.662414550781
    im_multiplicator(369) <= "1101000000001110"; --- j-0.749145507812
    re_multiplicator(370) <= "1100111110001010"; ---  -0.757202148438
    im_multiplicator(370) <= "1101011000110010"; --- j-0.653198242188
    re_multiplicator(371) <= "1100101001011011"; ---  -0.838195800781
    im_multiplicator(371) <= "1101110100011001"; --- j-0.545349121094
    re_multiplicator(372) <= "1100011000100101"; ---  -0.903991699219
    im_multiplicator(372) <= "1110010010100011"; --- j-0.427551269531
    re_multiplicator(373) <= "1100001011111101"; ---  -0.953308105469
    im_multiplicator(373) <= "1110110010101100"; --- j-0.302001953125
    re_multiplicator(374) <= "1100000011110001"; ---  -0.985290527344
    im_multiplicator(374) <= "1111010100001111"; --- j-0.170959472656
    re_multiplicator(375) <= "1100000000001011"; ---  -0.999328613281
    im_multiplicator(375) <= "1111110110100101"; --- j-0.0368041992188
    re_multiplicator(376) <= "1100000001001111"; ---  -0.995178222656
    im_multiplicator(376) <= "0000011001000110"; --- j0.0980224609375
    re_multiplicator(377) <= "1100000110111011"; ---  -0.972961425781
    im_multiplicator(377) <= "0000111011001010"; --- j0.231079101562
    re_multiplicator(378) <= "1100010001001010"; ---  -0.932983398438
    im_multiplicator(378) <= "0001011100001001"; --- j0.359924316406
    re_multiplicator(379) <= "1100011111101110"; ---  -0.876098632812
    im_multiplicator(379) <= "0001111011011100"; --- j0.482177734375
    re_multiplicator(380) <= "1100110010011000"; ---  -0.80322265625
    im_multiplicator(380) <= "0010011000100000"; --- j0.595703125
    re_multiplicator(381) <= "1101001000110001"; ---  -0.715759277344
    im_multiplicator(381) <= "0010110010110010"; --- j0.698364257812
    re_multiplicator(382) <= "1101100010100000"; ---  -0.615234375
    im_multiplicator(382) <= "0011001001110100"; --- j0.788330078125
    re_multiplicator(383) <= "1101111111000110"; ---  -0.503540039062
    im_multiplicator(383) <= "0011011101001011"; --- j0.863952636719
    re_multiplicator(385) <= "0011111101001111"; ---  0.989196777344
    im_multiplicator(385) <= "1111011010011100"; --- j-0.146728515625
    re_multiplicator(386) <= "0011110100111111"; ---  0.956970214844
    im_multiplicator(386) <= "1110110101101100"; --- j-0.290283203125
    re_multiplicator(387) <= "0011100111011011"; ---  0.903991699219
    im_multiplicator(387) <= "1110010010100011"; --- j-0.427551269531
    re_multiplicator(388) <= "0011010100110111"; ---  0.831481933594
    im_multiplicator(388) <= "1101110001110010"; --- j-0.555541992188
    re_multiplicator(389) <= "0010111101101100"; ---  0.740966796875
    im_multiplicator(389) <= "1101010100000101"; --- j-0.671569824219
    re_multiplicator(390) <= "0010100010011010"; ---  0.634399414062
    im_multiplicator(390) <= "1100111010000111"; --- j-0.773010253906
    re_multiplicator(391) <= "0010000011100111"; ---  0.514099121094
    im_multiplicator(391) <= "1100100100011011"; --- j-0.857727050781
    re_multiplicator(392) <= "0001100001111110"; ---  0.382690429688
    im_multiplicator(392) <= "1100010011011111"; --- j-0.923889160156
    re_multiplicator(393) <= "0000111110001101"; ---  0.242980957031
    im_multiplicator(393) <= "1100000111101011"; --- j-0.970031738281
    re_multiplicator(394) <= "0000011001000110"; ---  0.0980224609375
    im_multiplicator(394) <= "1100000001001111"; --- j-0.995178222656
    re_multiplicator(395) <= "1111110011011100"; ---  -0.049072265625
    im_multiplicator(395) <= "1100000000010100"; --- j-0.998779296875
    re_multiplicator(396) <= "1111001110000100"; ---  -0.195068359375
    im_multiplicator(396) <= "1100000100111011"; --- j-0.980773925781
    re_multiplicator(397) <= "1110101001110000"; ---  -0.3369140625
    im_multiplicator(397) <= "1100001110111110"; --- j-0.941528320312
    re_multiplicator(398) <= "1110000111010101"; ---  -0.471374511719
    im_multiplicator(398) <= "1100011110001111"; --- j-0.881896972656
    re_multiplicator(399) <= "1101100111100000"; ---  -0.595703125
    im_multiplicator(399) <= "1100110010011000"; --- j-0.80322265625
    re_multiplicator(400) <= "1101001010111111"; ---  -0.707092285156
    im_multiplicator(400) <= "1101001010111111"; --- j-0.707092285156
    re_multiplicator(401) <= "1100110010011000"; ---  -0.80322265625
    im_multiplicator(401) <= "1101100111100000"; --- j-0.595703125
    re_multiplicator(402) <= "1100011110001111"; ---  -0.881896972656
    im_multiplicator(402) <= "1110000111010101"; --- j-0.471374511719
    re_multiplicator(403) <= "1100001110111110"; ---  -0.941528320312
    im_multiplicator(403) <= "1110101001110000"; --- j-0.3369140625
    re_multiplicator(404) <= "1100000100111011"; ---  -0.980773925781
    im_multiplicator(404) <= "1111001110000100"; --- j-0.195068359375
    re_multiplicator(405) <= "1100000000010100"; ---  -0.998779296875
    im_multiplicator(405) <= "1111110011011100"; --- j-0.049072265625
    re_multiplicator(406) <= "1100000001001111"; ---  -0.995178222656
    im_multiplicator(406) <= "0000011001000110"; --- j0.0980224609375
    re_multiplicator(407) <= "1100000111101011"; ---  -0.970031738281
    im_multiplicator(407) <= "0000111110001101"; --- j0.242980957031
    re_multiplicator(408) <= "1100010011011111"; ---  -0.923889160156
    im_multiplicator(408) <= "0001100001111110"; --- j0.382690429688
    re_multiplicator(409) <= "1100100100011011"; ---  -0.857727050781
    im_multiplicator(409) <= "0010000011100111"; --- j0.514099121094
    re_multiplicator(410) <= "1100111010000111"; ---  -0.773010253906
    im_multiplicator(410) <= "0010100010011010"; --- j0.634399414062
    re_multiplicator(411) <= "1101010100000101"; ---  -0.671569824219
    im_multiplicator(411) <= "0010111101101100"; --- j0.740966796875
    re_multiplicator(412) <= "1101110001110010"; ---  -0.555541992188
    im_multiplicator(412) <= "0011010100110111"; --- j0.831481933594
    re_multiplicator(413) <= "1110010010100011"; ---  -0.427551269531
    im_multiplicator(413) <= "0011100111011011"; --- j0.903991699219
    re_multiplicator(414) <= "1110110101101100"; ---  -0.290283203125
    im_multiplicator(414) <= "0011110100111111"; --- j0.956970214844
    re_multiplicator(415) <= "1111011010011100"; ---  -0.146728515625
    im_multiplicator(415) <= "0011111101001111"; --- j0.989196777344
    re_multiplicator(417) <= "0011111100110000"; ---  0.9873046875
    im_multiplicator(417) <= "1111010111010101"; --- j-0.158874511719
    re_multiplicator(418) <= "0011110011000101"; ---  0.949523925781
    im_multiplicator(418) <= "1110101111101101"; --- j-0.313659667969
    re_multiplicator(419) <= "0011100011001111"; ---  0.887634277344
    im_multiplicator(419) <= "1110001010000111"; --- j-0.460510253906
    re_multiplicator(420) <= "0011001101101000"; ---  0.80322265625
    im_multiplicator(420) <= "1101100111100000"; --- j-0.595703125
    re_multiplicator(421) <= "0010110010110010"; ---  0.698364257812
    im_multiplicator(421) <= "1101001000110001"; --- j-0.715759277344
    re_multiplicator(422) <= "0010010011011010"; ---  0.575805664062
    im_multiplicator(422) <= "1100101110101101"; --- j-0.817565917969
    re_multiplicator(423) <= "0001110000010010"; ---  0.438598632812
    im_multiplicator(423) <= "1100011001111100"; --- j-0.898681640625
    re_multiplicator(424) <= "0001001010010100"; ---  0.290283203125
    im_multiplicator(424) <= "1100001011000001"; --- j-0.956970214844
    re_multiplicator(425) <= "0000100010011101"; ---  0.134582519531
    im_multiplicator(425) <= "1100000010010101"; --- j-0.990905761719
    re_multiplicator(426) <= "1111111001101110"; ---  -0.0245361328125
    im_multiplicator(426) <= "1100000000000101"; --- j-0.999694824219
    re_multiplicator(427) <= "1111010001001001"; ---  -0.183044433594
    im_multiplicator(427) <= "1100000100010101"; --- j-0.983093261719
    re_multiplicator(428) <= "1110101001110000"; ---  -0.3369140625
    im_multiplicator(428) <= "1100001110111110"; --- j-0.941528320312
    re_multiplicator(429) <= "1110000100100100"; ---  -0.482177734375
    im_multiplicator(429) <= "1100011111101110"; --- j-0.876098632812
    re_multiplicator(430) <= "1101100010100000"; ---  -0.615234375
    im_multiplicator(430) <= "1100110110001100"; --- j-0.788330078125
    re_multiplicator(431) <= "1101000100011100"; ---  -0.732666015625
    im_multiplicator(431) <= "1101010001110001"; --- j-0.680603027344
    re_multiplicator(432) <= "1100101011001001"; ---  -0.831481933594
    im_multiplicator(432) <= "1101110001110010"; --- j-0.555541992188
    re_multiplicator(433) <= "1100010111010000"; ---  -0.9091796875
    im_multiplicator(433) <= "1110010101011001"; --- j-0.416442871094
    re_multiplicator(434) <= "1100001001010001"; ---  -0.963806152344
    im_multiplicator(434) <= "1110111011101110"; --- j-0.266723632812
    re_multiplicator(435) <= "1100000001100100"; ---  -0.993896484375
    im_multiplicator(435) <= "1111100011110010"; --- j-0.110229492188
    re_multiplicator(436) <= "1100000000010100"; ---  -0.998779296875
    im_multiplicator(436) <= "0000001100100100"; --- j0.049072265625
    re_multiplicator(437) <= "1100000101100011"; ---  -0.978332519531
    im_multiplicator(437) <= "0000110101000001"; --- j0.207092285156
    re_multiplicator(438) <= "1100010001001010"; ---  -0.932983398438
    im_multiplicator(438) <= "0001011100001001"; --- j0.359924316406
    re_multiplicator(439) <= "1100100010110101"; ---  -0.863952636719
    im_multiplicator(439) <= "0010000000111010"; --- j0.503540039062
    re_multiplicator(440) <= "1100111010000111"; ---  -0.773010253906
    im_multiplicator(440) <= "0010100010011010"; --- j0.634399414062
    re_multiplicator(441) <= "1101010110011011"; ---  -0.662414550781
    im_multiplicator(441) <= "0010111111110010"; --- j0.749145507812
    re_multiplicator(442) <= "1101110111000011"; ---  -0.534973144531
    im_multiplicator(442) <= "0011011000010010"; --- j0.844848632812
    re_multiplicator(443) <= "1110011011001001"; ---  -0.393981933594
    im_multiplicator(443) <= "0011101011010011"; --- j0.919128417969
    re_multiplicator(444) <= "1111000001110011"; ---  -0.242980957031
    im_multiplicator(444) <= "0011111000010101"; --- j0.970031738281
    re_multiplicator(445) <= "1111101010000010"; ---  -0.0858154296875
    im_multiplicator(445) <= "0011111111000100"; --- j0.996337890625
    re_multiplicator(446) <= "0000010010110101"; ---  0.0735473632812
    im_multiplicator(446) <= "0011111111010100"; --- j0.997314453125
    re_multiplicator(447) <= "0000111011001010"; ---  0.231079101562
    im_multiplicator(447) <= "0011111001000101"; --- j0.972961425781
    re_multiplicator(449) <= "0011111100001111"; ---  0.985290527344
    im_multiplicator(449) <= "1111010100001111"; --- j-0.170959472656
    re_multiplicator(450) <= "0011110001000010"; ---  0.941528320312
    im_multiplicator(450) <= "1110101001110000"; --- j-0.3369140625
    re_multiplicator(451) <= "0011011110110000"; ---  0.8701171875
    im_multiplicator(451) <= "1110000001110100"; --- j-0.492919921875
    re_multiplicator(452) <= "0011000101111001"; ---  0.773010253906
    im_multiplicator(452) <= "1101011101100110"; --- j-0.634399414062
    re_multiplicator(453) <= "0010100111001110"; ---  0.653198242188
    im_multiplicator(453) <= "1100111110001010"; --- j-0.757202148438
    re_multiplicator(454) <= "0010000011100111"; ---  0.514099121094
    im_multiplicator(454) <= "1100100100011011"; --- j-0.857727050781
    re_multiplicator(455) <= "0001011100001001"; ---  0.359924316406
    im_multiplicator(455) <= "1100010001001010"; --- j-0.932983398438
    re_multiplicator(456) <= "0000110001111100"; ---  0.195068359375
    im_multiplicator(456) <= "1100000100111011"; --- j-0.980773925781
    re_multiplicator(457) <= "0000000110010010"; ---  0.0245361328125
    im_multiplicator(457) <= "1100000000000101"; --- j-0.999694824219
    re_multiplicator(458) <= "1111011010011100"; ---  -0.146728515625
    im_multiplicator(458) <= "1100000010110001"; --- j-0.989196777344
    re_multiplicator(459) <= "1110101111101101"; ---  -0.313659667969
    im_multiplicator(459) <= "1100001100111011"; --- j-0.949523925781
    re_multiplicator(460) <= "1110000111010101"; ---  -0.471374511719
    im_multiplicator(460) <= "1100011110001111"; --- j-0.881896972656
    re_multiplicator(461) <= "1101100010100000"; ---  -0.615234375
    im_multiplicator(461) <= "1100110110001100"; --- j-0.788330078125
    re_multiplicator(462) <= "1101000010010100"; ---  -0.740966796875
    im_multiplicator(462) <= "1101010100000101"; --- j-0.671569824219
    re_multiplicator(463) <= "1100100111101110"; ---  -0.844848632812
    im_multiplicator(463) <= "1101110111000011"; --- j-0.534973144531
    re_multiplicator(464) <= "1100010011011111"; ---  -0.923889160156
    im_multiplicator(464) <= "1110011110000010"; --- j-0.382690429688
    re_multiplicator(465) <= "1100000110001110"; ---  -0.975708007812
    im_multiplicator(465) <= "1111000111111010"; --- j-0.219116210938
    re_multiplicator(466) <= "1100000000010100"; ---  -0.998779296875
    im_multiplicator(466) <= "1111110011011100"; --- j-0.049072265625
    re_multiplicator(467) <= "1100000001111011"; ---  -0.992492675781
    im_multiplicator(467) <= "0000011111010110"; --- j0.122436523438
    re_multiplicator(468) <= "1100001011000001"; ---  -0.956970214844
    im_multiplicator(468) <= "0001001010010100"; --- j0.290283203125
    re_multiplicator(469) <= "1100011011010101"; ---  -0.893249511719
    im_multiplicator(469) <= "0001110011000110"; --- j0.449584960938
    re_multiplicator(470) <= "1100110010011000"; ---  -0.80322265625
    im_multiplicator(470) <= "0010011000100000"; --- j0.595703125
    re_multiplicator(471) <= "1101001111011111"; ---  -0.689514160156
    im_multiplicator(471) <= "0010111001011010"; --- j0.724243164062
    re_multiplicator(472) <= "1101110001110010"; ---  -0.555541992188
    im_multiplicator(472) <= "0011010100110111"; --- j0.831481933594
    re_multiplicator(473) <= "1110011000010001"; ---  -0.405212402344
    im_multiplicator(473) <= "0011101010000010"; --- j0.914184570312
    re_multiplicator(474) <= "1111000001110011"; ---  -0.242980957031
    im_multiplicator(474) <= "0011111000010101"; --- j0.970031738281
    re_multiplicator(475) <= "1111101101001011"; ---  -0.0735473632812
    im_multiplicator(475) <= "0011111111010100"; --- j0.997314453125
    re_multiplicator(476) <= "0000011001000110"; ---  0.0980224609375
    im_multiplicator(476) <= "0011111110110001"; --- j0.995178222656
    re_multiplicator(477) <= "0001000100010010"; ---  0.266723632812
    im_multiplicator(477) <= "0011110110101111"; --- j0.963806152344
    re_multiplicator(478) <= "0001101101011101"; ---  0.427551269531
    im_multiplicator(478) <= "0011100111011011"; --- j0.903991699219
    re_multiplicator(479) <= "0010010011011010"; ---  0.575805664062
    im_multiplicator(479) <= "0011010001010011"; --- j0.817565917969
    re_multiplicator(481) <= "0011111011101011"; ---  0.983093261719
    im_multiplicator(481) <= "1111010001001001"; --- j-0.183044433594
    re_multiplicator(482) <= "0011101110110110"; ---  0.932983398438
    im_multiplicator(482) <= "1110100011110111"; --- j-0.359924316406
    re_multiplicator(483) <= "0011011001111101"; ---  0.851379394531
    im_multiplicator(483) <= "1101111001101101"; --- j-0.524597167969
    re_multiplicator(484) <= "0010111101101100"; ---  0.740966796875
    im_multiplicator(484) <= "1101010100000101"; --- j-0.671569824219
    re_multiplicator(485) <= "0010011011000001"; ---  0.605529785156
    im_multiplicator(485) <= "1100110100010001"; --- j-0.795837402344
    re_multiplicator(486) <= "0001110011000110"; ---  0.449584960938
    im_multiplicator(486) <= "1100011011010101"; --- j-0.893249511719
    re_multiplicator(487) <= "0001000111010011"; ---  0.278503417969
    im_multiplicator(487) <= "1100001010001000"; --- j-0.96044921875
    re_multiplicator(488) <= "0000011001000110"; ---  0.0980224609375
    im_multiplicator(488) <= "1100000001001111"; --- j-0.995178222656
    re_multiplicator(489) <= "1111101010000010"; ---  -0.0858154296875
    im_multiplicator(489) <= "1100000000111100"; --- j-0.996337890625
    re_multiplicator(490) <= "1110111011101110"; ---  -0.266723632812
    im_multiplicator(490) <= "1100001001010001"; --- j-0.963806152344
    re_multiplicator(491) <= "1110001111101110"; ---  -0.438598632812
    im_multiplicator(491) <= "1100011001111100"; --- j-0.898681640625
    re_multiplicator(492) <= "1101100111100000"; ---  -0.595703125
    im_multiplicator(492) <= "1100110010011000"; --- j-0.80322265625
    re_multiplicator(493) <= "1101000100011100"; ---  -0.732666015625
    im_multiplicator(493) <= "1101010001110001"; --- j-0.680603027344
    re_multiplicator(494) <= "1100100111101110"; ---  -0.844848632812
    im_multiplicator(494) <= "1101110111000011"; --- j-0.534973144531
    re_multiplicator(495) <= "1100010010010011"; ---  -0.928527832031
    im_multiplicator(495) <= "1110100000111100"; --- j-0.371337890625
    re_multiplicator(496) <= "1100000100111011"; ---  -0.980773925781
    im_multiplicator(496) <= "1111001110000100"; --- j-0.195068359375
    re_multiplicator(497) <= "1100000000000001"; ---  -0.999938964844
    im_multiplicator(497) <= "1111111100110111"; --- j-0.0122680664062
    re_multiplicator(498) <= "1100000011110001"; ---  -0.985290527344
    im_multiplicator(498) <= "0000101011110001"; --- j0.170959472656
    re_multiplicator(499) <= "1100010000000011"; ---  -0.937316894531
    im_multiplicator(499) <= "0001011001001100"; --- j0.348388671875
    re_multiplicator(500) <= "1100100100011011"; ---  -0.857727050781
    im_multiplicator(500) <= "0010000011100111"; --- j0.514099121094
    re_multiplicator(501) <= "1101000000001110"; ---  -0.749145507812
    im_multiplicator(501) <= "0010101001100101"; --- j0.662414550781
    re_multiplicator(502) <= "1101100010100000"; ---  -0.615234375
    im_multiplicator(502) <= "0011001001110100"; --- j0.788330078125
    re_multiplicator(503) <= "1110001010000111"; ---  -0.460510253906
    im_multiplicator(503) <= "0011100011001111"; --- j0.887634277344
    re_multiplicator(504) <= "1110110101101100"; ---  -0.290283203125
    im_multiplicator(504) <= "0011110100111111"; --- j0.956970214844
    re_multiplicator(505) <= "1111100011110010"; ---  -0.110229492188
    im_multiplicator(505) <= "0011111110011100"; --- j0.993896484375
    re_multiplicator(506) <= "0000010010110101"; ---  0.0735473632812
    im_multiplicator(506) <= "0011111111010100"; --- j0.997314453125
    re_multiplicator(507) <= "0001000001010000"; ---  0.2548828125
    im_multiplicator(507) <= "0011110111100011"; --- j0.966979980469
    re_multiplicator(508) <= "0001101101011101"; ---  0.427551269531
    im_multiplicator(508) <= "0011100111011011"; --- j0.903991699219
    re_multiplicator(509) <= "0010010101111110"; ---  0.585815429688
    im_multiplicator(509) <= "0011001111011111"; --- j0.810485839844
    re_multiplicator(510) <= "0010111001011010"; ---  0.724243164062
    im_multiplicator(510) <= "0010110000100001"; --- j0.689514160156
    re_multiplicator(511) <= "0011010110100101"; ---  0.838195800781
    im_multiplicator(511) <= "0010001011100111"; --- j0.545349121094

    tmp_first_stage_re_out <= first_stage_re_out;
    tmp_first_stage_im_out <= first_stage_im_out;
    tmp_mul_re_out <= mul_re_out;
    tmp_mul_im_out <= mul_im_out;

    --- left-hand-side processors
    ULFFT_PT16_0 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(0),
            data_re_in(1) => data_re_in(32),
            data_re_in(2) => data_re_in(64),
            data_re_in(3) => data_re_in(96),
            data_re_in(4) => data_re_in(128),
            data_re_in(5) => data_re_in(160),
            data_re_in(6) => data_re_in(192),
            data_re_in(7) => data_re_in(224),
            data_re_in(8) => data_re_in(256),
            data_re_in(9) => data_re_in(288),
            data_re_in(10) => data_re_in(320),
            data_re_in(11) => data_re_in(352),
            data_re_in(12) => data_re_in(384),
            data_re_in(13) => data_re_in(416),
            data_re_in(14) => data_re_in(448),
            data_re_in(15) => data_re_in(480),
            data_im_in(0) => data_im_in(0),
            data_im_in(1) => data_im_in(32),
            data_im_in(2) => data_im_in(64),
            data_im_in(3) => data_im_in(96),
            data_im_in(4) => data_im_in(128),
            data_im_in(5) => data_im_in(160),
            data_im_in(6) => data_im_in(192),
            data_im_in(7) => data_im_in(224),
            data_im_in(8) => data_im_in(256),
            data_im_in(9) => data_im_in(288),
            data_im_in(10) => data_im_in(320),
            data_im_in(11) => data_im_in(352),
            data_im_in(12) => data_im_in(384),
            data_im_in(13) => data_im_in(416),
            data_im_in(14) => data_im_in(448),
            data_im_in(15) => data_im_in(480),
            data_re_out(0) => first_stage_re_out(0),
            data_re_out(1) => first_stage_re_out(32),
            data_re_out(2) => first_stage_re_out(64),
            data_re_out(3) => first_stage_re_out(96),
            data_re_out(4) => first_stage_re_out(128),
            data_re_out(5) => first_stage_re_out(160),
            data_re_out(6) => first_stage_re_out(192),
            data_re_out(7) => first_stage_re_out(224),
            data_re_out(8) => first_stage_re_out(256),
            data_re_out(9) => first_stage_re_out(288),
            data_re_out(10) => first_stage_re_out(320),
            data_re_out(11) => first_stage_re_out(352),
            data_re_out(12) => first_stage_re_out(384),
            data_re_out(13) => first_stage_re_out(416),
            data_re_out(14) => first_stage_re_out(448),
            data_re_out(15) => first_stage_re_out(480),
            data_im_out(0) => first_stage_im_out(0),
            data_im_out(1) => first_stage_im_out(32),
            data_im_out(2) => first_stage_im_out(64),
            data_im_out(3) => first_stage_im_out(96),
            data_im_out(4) => first_stage_im_out(128),
            data_im_out(5) => first_stage_im_out(160),
            data_im_out(6) => first_stage_im_out(192),
            data_im_out(7) => first_stage_im_out(224),
            data_im_out(8) => first_stage_im_out(256),
            data_im_out(9) => first_stage_im_out(288),
            data_im_out(10) => first_stage_im_out(320),
            data_im_out(11) => first_stage_im_out(352),
            data_im_out(12) => first_stage_im_out(384),
            data_im_out(13) => first_stage_im_out(416),
            data_im_out(14) => first_stage_im_out(448),
            data_im_out(15) => first_stage_im_out(480)
        );

    ULFFT_PT16_1 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(1),
            data_re_in(1) => data_re_in(33),
            data_re_in(2) => data_re_in(65),
            data_re_in(3) => data_re_in(97),
            data_re_in(4) => data_re_in(129),
            data_re_in(5) => data_re_in(161),
            data_re_in(6) => data_re_in(193),
            data_re_in(7) => data_re_in(225),
            data_re_in(8) => data_re_in(257),
            data_re_in(9) => data_re_in(289),
            data_re_in(10) => data_re_in(321),
            data_re_in(11) => data_re_in(353),
            data_re_in(12) => data_re_in(385),
            data_re_in(13) => data_re_in(417),
            data_re_in(14) => data_re_in(449),
            data_re_in(15) => data_re_in(481),
            data_im_in(0) => data_im_in(1),
            data_im_in(1) => data_im_in(33),
            data_im_in(2) => data_im_in(65),
            data_im_in(3) => data_im_in(97),
            data_im_in(4) => data_im_in(129),
            data_im_in(5) => data_im_in(161),
            data_im_in(6) => data_im_in(193),
            data_im_in(7) => data_im_in(225),
            data_im_in(8) => data_im_in(257),
            data_im_in(9) => data_im_in(289),
            data_im_in(10) => data_im_in(321),
            data_im_in(11) => data_im_in(353),
            data_im_in(12) => data_im_in(385),
            data_im_in(13) => data_im_in(417),
            data_im_in(14) => data_im_in(449),
            data_im_in(15) => data_im_in(481),
            data_re_out(0) => first_stage_re_out(1),
            data_re_out(1) => first_stage_re_out(33),
            data_re_out(2) => first_stage_re_out(65),
            data_re_out(3) => first_stage_re_out(97),
            data_re_out(4) => first_stage_re_out(129),
            data_re_out(5) => first_stage_re_out(161),
            data_re_out(6) => first_stage_re_out(193),
            data_re_out(7) => first_stage_re_out(225),
            data_re_out(8) => first_stage_re_out(257),
            data_re_out(9) => first_stage_re_out(289),
            data_re_out(10) => first_stage_re_out(321),
            data_re_out(11) => first_stage_re_out(353),
            data_re_out(12) => first_stage_re_out(385),
            data_re_out(13) => first_stage_re_out(417),
            data_re_out(14) => first_stage_re_out(449),
            data_re_out(15) => first_stage_re_out(481),
            data_im_out(0) => first_stage_im_out(1),
            data_im_out(1) => first_stage_im_out(33),
            data_im_out(2) => first_stage_im_out(65),
            data_im_out(3) => first_stage_im_out(97),
            data_im_out(4) => first_stage_im_out(129),
            data_im_out(5) => first_stage_im_out(161),
            data_im_out(6) => first_stage_im_out(193),
            data_im_out(7) => first_stage_im_out(225),
            data_im_out(8) => first_stage_im_out(257),
            data_im_out(9) => first_stage_im_out(289),
            data_im_out(10) => first_stage_im_out(321),
            data_im_out(11) => first_stage_im_out(353),
            data_im_out(12) => first_stage_im_out(385),
            data_im_out(13) => first_stage_im_out(417),
            data_im_out(14) => first_stage_im_out(449),
            data_im_out(15) => first_stage_im_out(481)
        );

    ULFFT_PT16_2 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(2),
            data_re_in(1) => data_re_in(34),
            data_re_in(2) => data_re_in(66),
            data_re_in(3) => data_re_in(98),
            data_re_in(4) => data_re_in(130),
            data_re_in(5) => data_re_in(162),
            data_re_in(6) => data_re_in(194),
            data_re_in(7) => data_re_in(226),
            data_re_in(8) => data_re_in(258),
            data_re_in(9) => data_re_in(290),
            data_re_in(10) => data_re_in(322),
            data_re_in(11) => data_re_in(354),
            data_re_in(12) => data_re_in(386),
            data_re_in(13) => data_re_in(418),
            data_re_in(14) => data_re_in(450),
            data_re_in(15) => data_re_in(482),
            data_im_in(0) => data_im_in(2),
            data_im_in(1) => data_im_in(34),
            data_im_in(2) => data_im_in(66),
            data_im_in(3) => data_im_in(98),
            data_im_in(4) => data_im_in(130),
            data_im_in(5) => data_im_in(162),
            data_im_in(6) => data_im_in(194),
            data_im_in(7) => data_im_in(226),
            data_im_in(8) => data_im_in(258),
            data_im_in(9) => data_im_in(290),
            data_im_in(10) => data_im_in(322),
            data_im_in(11) => data_im_in(354),
            data_im_in(12) => data_im_in(386),
            data_im_in(13) => data_im_in(418),
            data_im_in(14) => data_im_in(450),
            data_im_in(15) => data_im_in(482),
            data_re_out(0) => first_stage_re_out(2),
            data_re_out(1) => first_stage_re_out(34),
            data_re_out(2) => first_stage_re_out(66),
            data_re_out(3) => first_stage_re_out(98),
            data_re_out(4) => first_stage_re_out(130),
            data_re_out(5) => first_stage_re_out(162),
            data_re_out(6) => first_stage_re_out(194),
            data_re_out(7) => first_stage_re_out(226),
            data_re_out(8) => first_stage_re_out(258),
            data_re_out(9) => first_stage_re_out(290),
            data_re_out(10) => first_stage_re_out(322),
            data_re_out(11) => first_stage_re_out(354),
            data_re_out(12) => first_stage_re_out(386),
            data_re_out(13) => first_stage_re_out(418),
            data_re_out(14) => first_stage_re_out(450),
            data_re_out(15) => first_stage_re_out(482),
            data_im_out(0) => first_stage_im_out(2),
            data_im_out(1) => first_stage_im_out(34),
            data_im_out(2) => first_stage_im_out(66),
            data_im_out(3) => first_stage_im_out(98),
            data_im_out(4) => first_stage_im_out(130),
            data_im_out(5) => first_stage_im_out(162),
            data_im_out(6) => first_stage_im_out(194),
            data_im_out(7) => first_stage_im_out(226),
            data_im_out(8) => first_stage_im_out(258),
            data_im_out(9) => first_stage_im_out(290),
            data_im_out(10) => first_stage_im_out(322),
            data_im_out(11) => first_stage_im_out(354),
            data_im_out(12) => first_stage_im_out(386),
            data_im_out(13) => first_stage_im_out(418),
            data_im_out(14) => first_stage_im_out(450),
            data_im_out(15) => first_stage_im_out(482)
        );

    ULFFT_PT16_3 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(3),
            data_re_in(1) => data_re_in(35),
            data_re_in(2) => data_re_in(67),
            data_re_in(3) => data_re_in(99),
            data_re_in(4) => data_re_in(131),
            data_re_in(5) => data_re_in(163),
            data_re_in(6) => data_re_in(195),
            data_re_in(7) => data_re_in(227),
            data_re_in(8) => data_re_in(259),
            data_re_in(9) => data_re_in(291),
            data_re_in(10) => data_re_in(323),
            data_re_in(11) => data_re_in(355),
            data_re_in(12) => data_re_in(387),
            data_re_in(13) => data_re_in(419),
            data_re_in(14) => data_re_in(451),
            data_re_in(15) => data_re_in(483),
            data_im_in(0) => data_im_in(3),
            data_im_in(1) => data_im_in(35),
            data_im_in(2) => data_im_in(67),
            data_im_in(3) => data_im_in(99),
            data_im_in(4) => data_im_in(131),
            data_im_in(5) => data_im_in(163),
            data_im_in(6) => data_im_in(195),
            data_im_in(7) => data_im_in(227),
            data_im_in(8) => data_im_in(259),
            data_im_in(9) => data_im_in(291),
            data_im_in(10) => data_im_in(323),
            data_im_in(11) => data_im_in(355),
            data_im_in(12) => data_im_in(387),
            data_im_in(13) => data_im_in(419),
            data_im_in(14) => data_im_in(451),
            data_im_in(15) => data_im_in(483),
            data_re_out(0) => first_stage_re_out(3),
            data_re_out(1) => first_stage_re_out(35),
            data_re_out(2) => first_stage_re_out(67),
            data_re_out(3) => first_stage_re_out(99),
            data_re_out(4) => first_stage_re_out(131),
            data_re_out(5) => first_stage_re_out(163),
            data_re_out(6) => first_stage_re_out(195),
            data_re_out(7) => first_stage_re_out(227),
            data_re_out(8) => first_stage_re_out(259),
            data_re_out(9) => first_stage_re_out(291),
            data_re_out(10) => first_stage_re_out(323),
            data_re_out(11) => first_stage_re_out(355),
            data_re_out(12) => first_stage_re_out(387),
            data_re_out(13) => first_stage_re_out(419),
            data_re_out(14) => first_stage_re_out(451),
            data_re_out(15) => first_stage_re_out(483),
            data_im_out(0) => first_stage_im_out(3),
            data_im_out(1) => first_stage_im_out(35),
            data_im_out(2) => first_stage_im_out(67),
            data_im_out(3) => first_stage_im_out(99),
            data_im_out(4) => first_stage_im_out(131),
            data_im_out(5) => first_stage_im_out(163),
            data_im_out(6) => first_stage_im_out(195),
            data_im_out(7) => first_stage_im_out(227),
            data_im_out(8) => first_stage_im_out(259),
            data_im_out(9) => first_stage_im_out(291),
            data_im_out(10) => first_stage_im_out(323),
            data_im_out(11) => first_stage_im_out(355),
            data_im_out(12) => first_stage_im_out(387),
            data_im_out(13) => first_stage_im_out(419),
            data_im_out(14) => first_stage_im_out(451),
            data_im_out(15) => first_stage_im_out(483)
        );

    ULFFT_PT16_4 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(4),
            data_re_in(1) => data_re_in(36),
            data_re_in(2) => data_re_in(68),
            data_re_in(3) => data_re_in(100),
            data_re_in(4) => data_re_in(132),
            data_re_in(5) => data_re_in(164),
            data_re_in(6) => data_re_in(196),
            data_re_in(7) => data_re_in(228),
            data_re_in(8) => data_re_in(260),
            data_re_in(9) => data_re_in(292),
            data_re_in(10) => data_re_in(324),
            data_re_in(11) => data_re_in(356),
            data_re_in(12) => data_re_in(388),
            data_re_in(13) => data_re_in(420),
            data_re_in(14) => data_re_in(452),
            data_re_in(15) => data_re_in(484),
            data_im_in(0) => data_im_in(4),
            data_im_in(1) => data_im_in(36),
            data_im_in(2) => data_im_in(68),
            data_im_in(3) => data_im_in(100),
            data_im_in(4) => data_im_in(132),
            data_im_in(5) => data_im_in(164),
            data_im_in(6) => data_im_in(196),
            data_im_in(7) => data_im_in(228),
            data_im_in(8) => data_im_in(260),
            data_im_in(9) => data_im_in(292),
            data_im_in(10) => data_im_in(324),
            data_im_in(11) => data_im_in(356),
            data_im_in(12) => data_im_in(388),
            data_im_in(13) => data_im_in(420),
            data_im_in(14) => data_im_in(452),
            data_im_in(15) => data_im_in(484),
            data_re_out(0) => first_stage_re_out(4),
            data_re_out(1) => first_stage_re_out(36),
            data_re_out(2) => first_stage_re_out(68),
            data_re_out(3) => first_stage_re_out(100),
            data_re_out(4) => first_stage_re_out(132),
            data_re_out(5) => first_stage_re_out(164),
            data_re_out(6) => first_stage_re_out(196),
            data_re_out(7) => first_stage_re_out(228),
            data_re_out(8) => first_stage_re_out(260),
            data_re_out(9) => first_stage_re_out(292),
            data_re_out(10) => first_stage_re_out(324),
            data_re_out(11) => first_stage_re_out(356),
            data_re_out(12) => first_stage_re_out(388),
            data_re_out(13) => first_stage_re_out(420),
            data_re_out(14) => first_stage_re_out(452),
            data_re_out(15) => first_stage_re_out(484),
            data_im_out(0) => first_stage_im_out(4),
            data_im_out(1) => first_stage_im_out(36),
            data_im_out(2) => first_stage_im_out(68),
            data_im_out(3) => first_stage_im_out(100),
            data_im_out(4) => first_stage_im_out(132),
            data_im_out(5) => first_stage_im_out(164),
            data_im_out(6) => first_stage_im_out(196),
            data_im_out(7) => first_stage_im_out(228),
            data_im_out(8) => first_stage_im_out(260),
            data_im_out(9) => first_stage_im_out(292),
            data_im_out(10) => first_stage_im_out(324),
            data_im_out(11) => first_stage_im_out(356),
            data_im_out(12) => first_stage_im_out(388),
            data_im_out(13) => first_stage_im_out(420),
            data_im_out(14) => first_stage_im_out(452),
            data_im_out(15) => first_stage_im_out(484)
        );

    ULFFT_PT16_5 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(5),
            data_re_in(1) => data_re_in(37),
            data_re_in(2) => data_re_in(69),
            data_re_in(3) => data_re_in(101),
            data_re_in(4) => data_re_in(133),
            data_re_in(5) => data_re_in(165),
            data_re_in(6) => data_re_in(197),
            data_re_in(7) => data_re_in(229),
            data_re_in(8) => data_re_in(261),
            data_re_in(9) => data_re_in(293),
            data_re_in(10) => data_re_in(325),
            data_re_in(11) => data_re_in(357),
            data_re_in(12) => data_re_in(389),
            data_re_in(13) => data_re_in(421),
            data_re_in(14) => data_re_in(453),
            data_re_in(15) => data_re_in(485),
            data_im_in(0) => data_im_in(5),
            data_im_in(1) => data_im_in(37),
            data_im_in(2) => data_im_in(69),
            data_im_in(3) => data_im_in(101),
            data_im_in(4) => data_im_in(133),
            data_im_in(5) => data_im_in(165),
            data_im_in(6) => data_im_in(197),
            data_im_in(7) => data_im_in(229),
            data_im_in(8) => data_im_in(261),
            data_im_in(9) => data_im_in(293),
            data_im_in(10) => data_im_in(325),
            data_im_in(11) => data_im_in(357),
            data_im_in(12) => data_im_in(389),
            data_im_in(13) => data_im_in(421),
            data_im_in(14) => data_im_in(453),
            data_im_in(15) => data_im_in(485),
            data_re_out(0) => first_stage_re_out(5),
            data_re_out(1) => first_stage_re_out(37),
            data_re_out(2) => first_stage_re_out(69),
            data_re_out(3) => first_stage_re_out(101),
            data_re_out(4) => first_stage_re_out(133),
            data_re_out(5) => first_stage_re_out(165),
            data_re_out(6) => first_stage_re_out(197),
            data_re_out(7) => first_stage_re_out(229),
            data_re_out(8) => first_stage_re_out(261),
            data_re_out(9) => first_stage_re_out(293),
            data_re_out(10) => first_stage_re_out(325),
            data_re_out(11) => first_stage_re_out(357),
            data_re_out(12) => first_stage_re_out(389),
            data_re_out(13) => first_stage_re_out(421),
            data_re_out(14) => first_stage_re_out(453),
            data_re_out(15) => first_stage_re_out(485),
            data_im_out(0) => first_stage_im_out(5),
            data_im_out(1) => first_stage_im_out(37),
            data_im_out(2) => first_stage_im_out(69),
            data_im_out(3) => first_stage_im_out(101),
            data_im_out(4) => first_stage_im_out(133),
            data_im_out(5) => first_stage_im_out(165),
            data_im_out(6) => first_stage_im_out(197),
            data_im_out(7) => first_stage_im_out(229),
            data_im_out(8) => first_stage_im_out(261),
            data_im_out(9) => first_stage_im_out(293),
            data_im_out(10) => first_stage_im_out(325),
            data_im_out(11) => first_stage_im_out(357),
            data_im_out(12) => first_stage_im_out(389),
            data_im_out(13) => first_stage_im_out(421),
            data_im_out(14) => first_stage_im_out(453),
            data_im_out(15) => first_stage_im_out(485)
        );

    ULFFT_PT16_6 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(6),
            data_re_in(1) => data_re_in(38),
            data_re_in(2) => data_re_in(70),
            data_re_in(3) => data_re_in(102),
            data_re_in(4) => data_re_in(134),
            data_re_in(5) => data_re_in(166),
            data_re_in(6) => data_re_in(198),
            data_re_in(7) => data_re_in(230),
            data_re_in(8) => data_re_in(262),
            data_re_in(9) => data_re_in(294),
            data_re_in(10) => data_re_in(326),
            data_re_in(11) => data_re_in(358),
            data_re_in(12) => data_re_in(390),
            data_re_in(13) => data_re_in(422),
            data_re_in(14) => data_re_in(454),
            data_re_in(15) => data_re_in(486),
            data_im_in(0) => data_im_in(6),
            data_im_in(1) => data_im_in(38),
            data_im_in(2) => data_im_in(70),
            data_im_in(3) => data_im_in(102),
            data_im_in(4) => data_im_in(134),
            data_im_in(5) => data_im_in(166),
            data_im_in(6) => data_im_in(198),
            data_im_in(7) => data_im_in(230),
            data_im_in(8) => data_im_in(262),
            data_im_in(9) => data_im_in(294),
            data_im_in(10) => data_im_in(326),
            data_im_in(11) => data_im_in(358),
            data_im_in(12) => data_im_in(390),
            data_im_in(13) => data_im_in(422),
            data_im_in(14) => data_im_in(454),
            data_im_in(15) => data_im_in(486),
            data_re_out(0) => first_stage_re_out(6),
            data_re_out(1) => first_stage_re_out(38),
            data_re_out(2) => first_stage_re_out(70),
            data_re_out(3) => first_stage_re_out(102),
            data_re_out(4) => first_stage_re_out(134),
            data_re_out(5) => first_stage_re_out(166),
            data_re_out(6) => first_stage_re_out(198),
            data_re_out(7) => first_stage_re_out(230),
            data_re_out(8) => first_stage_re_out(262),
            data_re_out(9) => first_stage_re_out(294),
            data_re_out(10) => first_stage_re_out(326),
            data_re_out(11) => first_stage_re_out(358),
            data_re_out(12) => first_stage_re_out(390),
            data_re_out(13) => first_stage_re_out(422),
            data_re_out(14) => first_stage_re_out(454),
            data_re_out(15) => first_stage_re_out(486),
            data_im_out(0) => first_stage_im_out(6),
            data_im_out(1) => first_stage_im_out(38),
            data_im_out(2) => first_stage_im_out(70),
            data_im_out(3) => first_stage_im_out(102),
            data_im_out(4) => first_stage_im_out(134),
            data_im_out(5) => first_stage_im_out(166),
            data_im_out(6) => first_stage_im_out(198),
            data_im_out(7) => first_stage_im_out(230),
            data_im_out(8) => first_stage_im_out(262),
            data_im_out(9) => first_stage_im_out(294),
            data_im_out(10) => first_stage_im_out(326),
            data_im_out(11) => first_stage_im_out(358),
            data_im_out(12) => first_stage_im_out(390),
            data_im_out(13) => first_stage_im_out(422),
            data_im_out(14) => first_stage_im_out(454),
            data_im_out(15) => first_stage_im_out(486)
        );

    ULFFT_PT16_7 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(7),
            data_re_in(1) => data_re_in(39),
            data_re_in(2) => data_re_in(71),
            data_re_in(3) => data_re_in(103),
            data_re_in(4) => data_re_in(135),
            data_re_in(5) => data_re_in(167),
            data_re_in(6) => data_re_in(199),
            data_re_in(7) => data_re_in(231),
            data_re_in(8) => data_re_in(263),
            data_re_in(9) => data_re_in(295),
            data_re_in(10) => data_re_in(327),
            data_re_in(11) => data_re_in(359),
            data_re_in(12) => data_re_in(391),
            data_re_in(13) => data_re_in(423),
            data_re_in(14) => data_re_in(455),
            data_re_in(15) => data_re_in(487),
            data_im_in(0) => data_im_in(7),
            data_im_in(1) => data_im_in(39),
            data_im_in(2) => data_im_in(71),
            data_im_in(3) => data_im_in(103),
            data_im_in(4) => data_im_in(135),
            data_im_in(5) => data_im_in(167),
            data_im_in(6) => data_im_in(199),
            data_im_in(7) => data_im_in(231),
            data_im_in(8) => data_im_in(263),
            data_im_in(9) => data_im_in(295),
            data_im_in(10) => data_im_in(327),
            data_im_in(11) => data_im_in(359),
            data_im_in(12) => data_im_in(391),
            data_im_in(13) => data_im_in(423),
            data_im_in(14) => data_im_in(455),
            data_im_in(15) => data_im_in(487),
            data_re_out(0) => first_stage_re_out(7),
            data_re_out(1) => first_stage_re_out(39),
            data_re_out(2) => first_stage_re_out(71),
            data_re_out(3) => first_stage_re_out(103),
            data_re_out(4) => first_stage_re_out(135),
            data_re_out(5) => first_stage_re_out(167),
            data_re_out(6) => first_stage_re_out(199),
            data_re_out(7) => first_stage_re_out(231),
            data_re_out(8) => first_stage_re_out(263),
            data_re_out(9) => first_stage_re_out(295),
            data_re_out(10) => first_stage_re_out(327),
            data_re_out(11) => first_stage_re_out(359),
            data_re_out(12) => first_stage_re_out(391),
            data_re_out(13) => first_stage_re_out(423),
            data_re_out(14) => first_stage_re_out(455),
            data_re_out(15) => first_stage_re_out(487),
            data_im_out(0) => first_stage_im_out(7),
            data_im_out(1) => first_stage_im_out(39),
            data_im_out(2) => first_stage_im_out(71),
            data_im_out(3) => first_stage_im_out(103),
            data_im_out(4) => first_stage_im_out(135),
            data_im_out(5) => first_stage_im_out(167),
            data_im_out(6) => first_stage_im_out(199),
            data_im_out(7) => first_stage_im_out(231),
            data_im_out(8) => first_stage_im_out(263),
            data_im_out(9) => first_stage_im_out(295),
            data_im_out(10) => first_stage_im_out(327),
            data_im_out(11) => first_stage_im_out(359),
            data_im_out(12) => first_stage_im_out(391),
            data_im_out(13) => first_stage_im_out(423),
            data_im_out(14) => first_stage_im_out(455),
            data_im_out(15) => first_stage_im_out(487)
        );

    ULFFT_PT16_8 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(8),
            data_re_in(1) => data_re_in(40),
            data_re_in(2) => data_re_in(72),
            data_re_in(3) => data_re_in(104),
            data_re_in(4) => data_re_in(136),
            data_re_in(5) => data_re_in(168),
            data_re_in(6) => data_re_in(200),
            data_re_in(7) => data_re_in(232),
            data_re_in(8) => data_re_in(264),
            data_re_in(9) => data_re_in(296),
            data_re_in(10) => data_re_in(328),
            data_re_in(11) => data_re_in(360),
            data_re_in(12) => data_re_in(392),
            data_re_in(13) => data_re_in(424),
            data_re_in(14) => data_re_in(456),
            data_re_in(15) => data_re_in(488),
            data_im_in(0) => data_im_in(8),
            data_im_in(1) => data_im_in(40),
            data_im_in(2) => data_im_in(72),
            data_im_in(3) => data_im_in(104),
            data_im_in(4) => data_im_in(136),
            data_im_in(5) => data_im_in(168),
            data_im_in(6) => data_im_in(200),
            data_im_in(7) => data_im_in(232),
            data_im_in(8) => data_im_in(264),
            data_im_in(9) => data_im_in(296),
            data_im_in(10) => data_im_in(328),
            data_im_in(11) => data_im_in(360),
            data_im_in(12) => data_im_in(392),
            data_im_in(13) => data_im_in(424),
            data_im_in(14) => data_im_in(456),
            data_im_in(15) => data_im_in(488),
            data_re_out(0) => first_stage_re_out(8),
            data_re_out(1) => first_stage_re_out(40),
            data_re_out(2) => first_stage_re_out(72),
            data_re_out(3) => first_stage_re_out(104),
            data_re_out(4) => first_stage_re_out(136),
            data_re_out(5) => first_stage_re_out(168),
            data_re_out(6) => first_stage_re_out(200),
            data_re_out(7) => first_stage_re_out(232),
            data_re_out(8) => first_stage_re_out(264),
            data_re_out(9) => first_stage_re_out(296),
            data_re_out(10) => first_stage_re_out(328),
            data_re_out(11) => first_stage_re_out(360),
            data_re_out(12) => first_stage_re_out(392),
            data_re_out(13) => first_stage_re_out(424),
            data_re_out(14) => first_stage_re_out(456),
            data_re_out(15) => first_stage_re_out(488),
            data_im_out(0) => first_stage_im_out(8),
            data_im_out(1) => first_stage_im_out(40),
            data_im_out(2) => first_stage_im_out(72),
            data_im_out(3) => first_stage_im_out(104),
            data_im_out(4) => first_stage_im_out(136),
            data_im_out(5) => first_stage_im_out(168),
            data_im_out(6) => first_stage_im_out(200),
            data_im_out(7) => first_stage_im_out(232),
            data_im_out(8) => first_stage_im_out(264),
            data_im_out(9) => first_stage_im_out(296),
            data_im_out(10) => first_stage_im_out(328),
            data_im_out(11) => first_stage_im_out(360),
            data_im_out(12) => first_stage_im_out(392),
            data_im_out(13) => first_stage_im_out(424),
            data_im_out(14) => first_stage_im_out(456),
            data_im_out(15) => first_stage_im_out(488)
        );

    ULFFT_PT16_9 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(9),
            data_re_in(1) => data_re_in(41),
            data_re_in(2) => data_re_in(73),
            data_re_in(3) => data_re_in(105),
            data_re_in(4) => data_re_in(137),
            data_re_in(5) => data_re_in(169),
            data_re_in(6) => data_re_in(201),
            data_re_in(7) => data_re_in(233),
            data_re_in(8) => data_re_in(265),
            data_re_in(9) => data_re_in(297),
            data_re_in(10) => data_re_in(329),
            data_re_in(11) => data_re_in(361),
            data_re_in(12) => data_re_in(393),
            data_re_in(13) => data_re_in(425),
            data_re_in(14) => data_re_in(457),
            data_re_in(15) => data_re_in(489),
            data_im_in(0) => data_im_in(9),
            data_im_in(1) => data_im_in(41),
            data_im_in(2) => data_im_in(73),
            data_im_in(3) => data_im_in(105),
            data_im_in(4) => data_im_in(137),
            data_im_in(5) => data_im_in(169),
            data_im_in(6) => data_im_in(201),
            data_im_in(7) => data_im_in(233),
            data_im_in(8) => data_im_in(265),
            data_im_in(9) => data_im_in(297),
            data_im_in(10) => data_im_in(329),
            data_im_in(11) => data_im_in(361),
            data_im_in(12) => data_im_in(393),
            data_im_in(13) => data_im_in(425),
            data_im_in(14) => data_im_in(457),
            data_im_in(15) => data_im_in(489),
            data_re_out(0) => first_stage_re_out(9),
            data_re_out(1) => first_stage_re_out(41),
            data_re_out(2) => first_stage_re_out(73),
            data_re_out(3) => first_stage_re_out(105),
            data_re_out(4) => first_stage_re_out(137),
            data_re_out(5) => first_stage_re_out(169),
            data_re_out(6) => first_stage_re_out(201),
            data_re_out(7) => first_stage_re_out(233),
            data_re_out(8) => first_stage_re_out(265),
            data_re_out(9) => first_stage_re_out(297),
            data_re_out(10) => first_stage_re_out(329),
            data_re_out(11) => first_stage_re_out(361),
            data_re_out(12) => first_stage_re_out(393),
            data_re_out(13) => first_stage_re_out(425),
            data_re_out(14) => first_stage_re_out(457),
            data_re_out(15) => first_stage_re_out(489),
            data_im_out(0) => first_stage_im_out(9),
            data_im_out(1) => first_stage_im_out(41),
            data_im_out(2) => first_stage_im_out(73),
            data_im_out(3) => first_stage_im_out(105),
            data_im_out(4) => first_stage_im_out(137),
            data_im_out(5) => first_stage_im_out(169),
            data_im_out(6) => first_stage_im_out(201),
            data_im_out(7) => first_stage_im_out(233),
            data_im_out(8) => first_stage_im_out(265),
            data_im_out(9) => first_stage_im_out(297),
            data_im_out(10) => first_stage_im_out(329),
            data_im_out(11) => first_stage_im_out(361),
            data_im_out(12) => first_stage_im_out(393),
            data_im_out(13) => first_stage_im_out(425),
            data_im_out(14) => first_stage_im_out(457),
            data_im_out(15) => first_stage_im_out(489)
        );

    ULFFT_PT16_10 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(10),
            data_re_in(1) => data_re_in(42),
            data_re_in(2) => data_re_in(74),
            data_re_in(3) => data_re_in(106),
            data_re_in(4) => data_re_in(138),
            data_re_in(5) => data_re_in(170),
            data_re_in(6) => data_re_in(202),
            data_re_in(7) => data_re_in(234),
            data_re_in(8) => data_re_in(266),
            data_re_in(9) => data_re_in(298),
            data_re_in(10) => data_re_in(330),
            data_re_in(11) => data_re_in(362),
            data_re_in(12) => data_re_in(394),
            data_re_in(13) => data_re_in(426),
            data_re_in(14) => data_re_in(458),
            data_re_in(15) => data_re_in(490),
            data_im_in(0) => data_im_in(10),
            data_im_in(1) => data_im_in(42),
            data_im_in(2) => data_im_in(74),
            data_im_in(3) => data_im_in(106),
            data_im_in(4) => data_im_in(138),
            data_im_in(5) => data_im_in(170),
            data_im_in(6) => data_im_in(202),
            data_im_in(7) => data_im_in(234),
            data_im_in(8) => data_im_in(266),
            data_im_in(9) => data_im_in(298),
            data_im_in(10) => data_im_in(330),
            data_im_in(11) => data_im_in(362),
            data_im_in(12) => data_im_in(394),
            data_im_in(13) => data_im_in(426),
            data_im_in(14) => data_im_in(458),
            data_im_in(15) => data_im_in(490),
            data_re_out(0) => first_stage_re_out(10),
            data_re_out(1) => first_stage_re_out(42),
            data_re_out(2) => first_stage_re_out(74),
            data_re_out(3) => first_stage_re_out(106),
            data_re_out(4) => first_stage_re_out(138),
            data_re_out(5) => first_stage_re_out(170),
            data_re_out(6) => first_stage_re_out(202),
            data_re_out(7) => first_stage_re_out(234),
            data_re_out(8) => first_stage_re_out(266),
            data_re_out(9) => first_stage_re_out(298),
            data_re_out(10) => first_stage_re_out(330),
            data_re_out(11) => first_stage_re_out(362),
            data_re_out(12) => first_stage_re_out(394),
            data_re_out(13) => first_stage_re_out(426),
            data_re_out(14) => first_stage_re_out(458),
            data_re_out(15) => first_stage_re_out(490),
            data_im_out(0) => first_stage_im_out(10),
            data_im_out(1) => first_stage_im_out(42),
            data_im_out(2) => first_stage_im_out(74),
            data_im_out(3) => first_stage_im_out(106),
            data_im_out(4) => first_stage_im_out(138),
            data_im_out(5) => first_stage_im_out(170),
            data_im_out(6) => first_stage_im_out(202),
            data_im_out(7) => first_stage_im_out(234),
            data_im_out(8) => first_stage_im_out(266),
            data_im_out(9) => first_stage_im_out(298),
            data_im_out(10) => first_stage_im_out(330),
            data_im_out(11) => first_stage_im_out(362),
            data_im_out(12) => first_stage_im_out(394),
            data_im_out(13) => first_stage_im_out(426),
            data_im_out(14) => first_stage_im_out(458),
            data_im_out(15) => first_stage_im_out(490)
        );

    ULFFT_PT16_11 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(11),
            data_re_in(1) => data_re_in(43),
            data_re_in(2) => data_re_in(75),
            data_re_in(3) => data_re_in(107),
            data_re_in(4) => data_re_in(139),
            data_re_in(5) => data_re_in(171),
            data_re_in(6) => data_re_in(203),
            data_re_in(7) => data_re_in(235),
            data_re_in(8) => data_re_in(267),
            data_re_in(9) => data_re_in(299),
            data_re_in(10) => data_re_in(331),
            data_re_in(11) => data_re_in(363),
            data_re_in(12) => data_re_in(395),
            data_re_in(13) => data_re_in(427),
            data_re_in(14) => data_re_in(459),
            data_re_in(15) => data_re_in(491),
            data_im_in(0) => data_im_in(11),
            data_im_in(1) => data_im_in(43),
            data_im_in(2) => data_im_in(75),
            data_im_in(3) => data_im_in(107),
            data_im_in(4) => data_im_in(139),
            data_im_in(5) => data_im_in(171),
            data_im_in(6) => data_im_in(203),
            data_im_in(7) => data_im_in(235),
            data_im_in(8) => data_im_in(267),
            data_im_in(9) => data_im_in(299),
            data_im_in(10) => data_im_in(331),
            data_im_in(11) => data_im_in(363),
            data_im_in(12) => data_im_in(395),
            data_im_in(13) => data_im_in(427),
            data_im_in(14) => data_im_in(459),
            data_im_in(15) => data_im_in(491),
            data_re_out(0) => first_stage_re_out(11),
            data_re_out(1) => first_stage_re_out(43),
            data_re_out(2) => first_stage_re_out(75),
            data_re_out(3) => first_stage_re_out(107),
            data_re_out(4) => first_stage_re_out(139),
            data_re_out(5) => first_stage_re_out(171),
            data_re_out(6) => first_stage_re_out(203),
            data_re_out(7) => first_stage_re_out(235),
            data_re_out(8) => first_stage_re_out(267),
            data_re_out(9) => first_stage_re_out(299),
            data_re_out(10) => first_stage_re_out(331),
            data_re_out(11) => first_stage_re_out(363),
            data_re_out(12) => first_stage_re_out(395),
            data_re_out(13) => first_stage_re_out(427),
            data_re_out(14) => first_stage_re_out(459),
            data_re_out(15) => first_stage_re_out(491),
            data_im_out(0) => first_stage_im_out(11),
            data_im_out(1) => first_stage_im_out(43),
            data_im_out(2) => first_stage_im_out(75),
            data_im_out(3) => first_stage_im_out(107),
            data_im_out(4) => first_stage_im_out(139),
            data_im_out(5) => first_stage_im_out(171),
            data_im_out(6) => first_stage_im_out(203),
            data_im_out(7) => first_stage_im_out(235),
            data_im_out(8) => first_stage_im_out(267),
            data_im_out(9) => first_stage_im_out(299),
            data_im_out(10) => first_stage_im_out(331),
            data_im_out(11) => first_stage_im_out(363),
            data_im_out(12) => first_stage_im_out(395),
            data_im_out(13) => first_stage_im_out(427),
            data_im_out(14) => first_stage_im_out(459),
            data_im_out(15) => first_stage_im_out(491)
        );

    ULFFT_PT16_12 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(12),
            data_re_in(1) => data_re_in(44),
            data_re_in(2) => data_re_in(76),
            data_re_in(3) => data_re_in(108),
            data_re_in(4) => data_re_in(140),
            data_re_in(5) => data_re_in(172),
            data_re_in(6) => data_re_in(204),
            data_re_in(7) => data_re_in(236),
            data_re_in(8) => data_re_in(268),
            data_re_in(9) => data_re_in(300),
            data_re_in(10) => data_re_in(332),
            data_re_in(11) => data_re_in(364),
            data_re_in(12) => data_re_in(396),
            data_re_in(13) => data_re_in(428),
            data_re_in(14) => data_re_in(460),
            data_re_in(15) => data_re_in(492),
            data_im_in(0) => data_im_in(12),
            data_im_in(1) => data_im_in(44),
            data_im_in(2) => data_im_in(76),
            data_im_in(3) => data_im_in(108),
            data_im_in(4) => data_im_in(140),
            data_im_in(5) => data_im_in(172),
            data_im_in(6) => data_im_in(204),
            data_im_in(7) => data_im_in(236),
            data_im_in(8) => data_im_in(268),
            data_im_in(9) => data_im_in(300),
            data_im_in(10) => data_im_in(332),
            data_im_in(11) => data_im_in(364),
            data_im_in(12) => data_im_in(396),
            data_im_in(13) => data_im_in(428),
            data_im_in(14) => data_im_in(460),
            data_im_in(15) => data_im_in(492),
            data_re_out(0) => first_stage_re_out(12),
            data_re_out(1) => first_stage_re_out(44),
            data_re_out(2) => first_stage_re_out(76),
            data_re_out(3) => first_stage_re_out(108),
            data_re_out(4) => first_stage_re_out(140),
            data_re_out(5) => first_stage_re_out(172),
            data_re_out(6) => first_stage_re_out(204),
            data_re_out(7) => first_stage_re_out(236),
            data_re_out(8) => first_stage_re_out(268),
            data_re_out(9) => first_stage_re_out(300),
            data_re_out(10) => first_stage_re_out(332),
            data_re_out(11) => first_stage_re_out(364),
            data_re_out(12) => first_stage_re_out(396),
            data_re_out(13) => first_stage_re_out(428),
            data_re_out(14) => first_stage_re_out(460),
            data_re_out(15) => first_stage_re_out(492),
            data_im_out(0) => first_stage_im_out(12),
            data_im_out(1) => first_stage_im_out(44),
            data_im_out(2) => first_stage_im_out(76),
            data_im_out(3) => first_stage_im_out(108),
            data_im_out(4) => first_stage_im_out(140),
            data_im_out(5) => first_stage_im_out(172),
            data_im_out(6) => first_stage_im_out(204),
            data_im_out(7) => first_stage_im_out(236),
            data_im_out(8) => first_stage_im_out(268),
            data_im_out(9) => first_stage_im_out(300),
            data_im_out(10) => first_stage_im_out(332),
            data_im_out(11) => first_stage_im_out(364),
            data_im_out(12) => first_stage_im_out(396),
            data_im_out(13) => first_stage_im_out(428),
            data_im_out(14) => first_stage_im_out(460),
            data_im_out(15) => first_stage_im_out(492)
        );

    ULFFT_PT16_13 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(13),
            data_re_in(1) => data_re_in(45),
            data_re_in(2) => data_re_in(77),
            data_re_in(3) => data_re_in(109),
            data_re_in(4) => data_re_in(141),
            data_re_in(5) => data_re_in(173),
            data_re_in(6) => data_re_in(205),
            data_re_in(7) => data_re_in(237),
            data_re_in(8) => data_re_in(269),
            data_re_in(9) => data_re_in(301),
            data_re_in(10) => data_re_in(333),
            data_re_in(11) => data_re_in(365),
            data_re_in(12) => data_re_in(397),
            data_re_in(13) => data_re_in(429),
            data_re_in(14) => data_re_in(461),
            data_re_in(15) => data_re_in(493),
            data_im_in(0) => data_im_in(13),
            data_im_in(1) => data_im_in(45),
            data_im_in(2) => data_im_in(77),
            data_im_in(3) => data_im_in(109),
            data_im_in(4) => data_im_in(141),
            data_im_in(5) => data_im_in(173),
            data_im_in(6) => data_im_in(205),
            data_im_in(7) => data_im_in(237),
            data_im_in(8) => data_im_in(269),
            data_im_in(9) => data_im_in(301),
            data_im_in(10) => data_im_in(333),
            data_im_in(11) => data_im_in(365),
            data_im_in(12) => data_im_in(397),
            data_im_in(13) => data_im_in(429),
            data_im_in(14) => data_im_in(461),
            data_im_in(15) => data_im_in(493),
            data_re_out(0) => first_stage_re_out(13),
            data_re_out(1) => first_stage_re_out(45),
            data_re_out(2) => first_stage_re_out(77),
            data_re_out(3) => first_stage_re_out(109),
            data_re_out(4) => first_stage_re_out(141),
            data_re_out(5) => first_stage_re_out(173),
            data_re_out(6) => first_stage_re_out(205),
            data_re_out(7) => first_stage_re_out(237),
            data_re_out(8) => first_stage_re_out(269),
            data_re_out(9) => first_stage_re_out(301),
            data_re_out(10) => first_stage_re_out(333),
            data_re_out(11) => first_stage_re_out(365),
            data_re_out(12) => first_stage_re_out(397),
            data_re_out(13) => first_stage_re_out(429),
            data_re_out(14) => first_stage_re_out(461),
            data_re_out(15) => first_stage_re_out(493),
            data_im_out(0) => first_stage_im_out(13),
            data_im_out(1) => first_stage_im_out(45),
            data_im_out(2) => first_stage_im_out(77),
            data_im_out(3) => first_stage_im_out(109),
            data_im_out(4) => first_stage_im_out(141),
            data_im_out(5) => first_stage_im_out(173),
            data_im_out(6) => first_stage_im_out(205),
            data_im_out(7) => first_stage_im_out(237),
            data_im_out(8) => first_stage_im_out(269),
            data_im_out(9) => first_stage_im_out(301),
            data_im_out(10) => first_stage_im_out(333),
            data_im_out(11) => first_stage_im_out(365),
            data_im_out(12) => first_stage_im_out(397),
            data_im_out(13) => first_stage_im_out(429),
            data_im_out(14) => first_stage_im_out(461),
            data_im_out(15) => first_stage_im_out(493)
        );

    ULFFT_PT16_14 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(14),
            data_re_in(1) => data_re_in(46),
            data_re_in(2) => data_re_in(78),
            data_re_in(3) => data_re_in(110),
            data_re_in(4) => data_re_in(142),
            data_re_in(5) => data_re_in(174),
            data_re_in(6) => data_re_in(206),
            data_re_in(7) => data_re_in(238),
            data_re_in(8) => data_re_in(270),
            data_re_in(9) => data_re_in(302),
            data_re_in(10) => data_re_in(334),
            data_re_in(11) => data_re_in(366),
            data_re_in(12) => data_re_in(398),
            data_re_in(13) => data_re_in(430),
            data_re_in(14) => data_re_in(462),
            data_re_in(15) => data_re_in(494),
            data_im_in(0) => data_im_in(14),
            data_im_in(1) => data_im_in(46),
            data_im_in(2) => data_im_in(78),
            data_im_in(3) => data_im_in(110),
            data_im_in(4) => data_im_in(142),
            data_im_in(5) => data_im_in(174),
            data_im_in(6) => data_im_in(206),
            data_im_in(7) => data_im_in(238),
            data_im_in(8) => data_im_in(270),
            data_im_in(9) => data_im_in(302),
            data_im_in(10) => data_im_in(334),
            data_im_in(11) => data_im_in(366),
            data_im_in(12) => data_im_in(398),
            data_im_in(13) => data_im_in(430),
            data_im_in(14) => data_im_in(462),
            data_im_in(15) => data_im_in(494),
            data_re_out(0) => first_stage_re_out(14),
            data_re_out(1) => first_stage_re_out(46),
            data_re_out(2) => first_stage_re_out(78),
            data_re_out(3) => first_stage_re_out(110),
            data_re_out(4) => first_stage_re_out(142),
            data_re_out(5) => first_stage_re_out(174),
            data_re_out(6) => first_stage_re_out(206),
            data_re_out(7) => first_stage_re_out(238),
            data_re_out(8) => first_stage_re_out(270),
            data_re_out(9) => first_stage_re_out(302),
            data_re_out(10) => first_stage_re_out(334),
            data_re_out(11) => first_stage_re_out(366),
            data_re_out(12) => first_stage_re_out(398),
            data_re_out(13) => first_stage_re_out(430),
            data_re_out(14) => first_stage_re_out(462),
            data_re_out(15) => first_stage_re_out(494),
            data_im_out(0) => first_stage_im_out(14),
            data_im_out(1) => first_stage_im_out(46),
            data_im_out(2) => first_stage_im_out(78),
            data_im_out(3) => first_stage_im_out(110),
            data_im_out(4) => first_stage_im_out(142),
            data_im_out(5) => first_stage_im_out(174),
            data_im_out(6) => first_stage_im_out(206),
            data_im_out(7) => first_stage_im_out(238),
            data_im_out(8) => first_stage_im_out(270),
            data_im_out(9) => first_stage_im_out(302),
            data_im_out(10) => first_stage_im_out(334),
            data_im_out(11) => first_stage_im_out(366),
            data_im_out(12) => first_stage_im_out(398),
            data_im_out(13) => first_stage_im_out(430),
            data_im_out(14) => first_stage_im_out(462),
            data_im_out(15) => first_stage_im_out(494)
        );

    ULFFT_PT16_15 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(15),
            data_re_in(1) => data_re_in(47),
            data_re_in(2) => data_re_in(79),
            data_re_in(3) => data_re_in(111),
            data_re_in(4) => data_re_in(143),
            data_re_in(5) => data_re_in(175),
            data_re_in(6) => data_re_in(207),
            data_re_in(7) => data_re_in(239),
            data_re_in(8) => data_re_in(271),
            data_re_in(9) => data_re_in(303),
            data_re_in(10) => data_re_in(335),
            data_re_in(11) => data_re_in(367),
            data_re_in(12) => data_re_in(399),
            data_re_in(13) => data_re_in(431),
            data_re_in(14) => data_re_in(463),
            data_re_in(15) => data_re_in(495),
            data_im_in(0) => data_im_in(15),
            data_im_in(1) => data_im_in(47),
            data_im_in(2) => data_im_in(79),
            data_im_in(3) => data_im_in(111),
            data_im_in(4) => data_im_in(143),
            data_im_in(5) => data_im_in(175),
            data_im_in(6) => data_im_in(207),
            data_im_in(7) => data_im_in(239),
            data_im_in(8) => data_im_in(271),
            data_im_in(9) => data_im_in(303),
            data_im_in(10) => data_im_in(335),
            data_im_in(11) => data_im_in(367),
            data_im_in(12) => data_im_in(399),
            data_im_in(13) => data_im_in(431),
            data_im_in(14) => data_im_in(463),
            data_im_in(15) => data_im_in(495),
            data_re_out(0) => first_stage_re_out(15),
            data_re_out(1) => first_stage_re_out(47),
            data_re_out(2) => first_stage_re_out(79),
            data_re_out(3) => first_stage_re_out(111),
            data_re_out(4) => first_stage_re_out(143),
            data_re_out(5) => first_stage_re_out(175),
            data_re_out(6) => first_stage_re_out(207),
            data_re_out(7) => first_stage_re_out(239),
            data_re_out(8) => first_stage_re_out(271),
            data_re_out(9) => first_stage_re_out(303),
            data_re_out(10) => first_stage_re_out(335),
            data_re_out(11) => first_stage_re_out(367),
            data_re_out(12) => first_stage_re_out(399),
            data_re_out(13) => first_stage_re_out(431),
            data_re_out(14) => first_stage_re_out(463),
            data_re_out(15) => first_stage_re_out(495),
            data_im_out(0) => first_stage_im_out(15),
            data_im_out(1) => first_stage_im_out(47),
            data_im_out(2) => first_stage_im_out(79),
            data_im_out(3) => first_stage_im_out(111),
            data_im_out(4) => first_stage_im_out(143),
            data_im_out(5) => first_stage_im_out(175),
            data_im_out(6) => first_stage_im_out(207),
            data_im_out(7) => first_stage_im_out(239),
            data_im_out(8) => first_stage_im_out(271),
            data_im_out(9) => first_stage_im_out(303),
            data_im_out(10) => first_stage_im_out(335),
            data_im_out(11) => first_stage_im_out(367),
            data_im_out(12) => first_stage_im_out(399),
            data_im_out(13) => first_stage_im_out(431),
            data_im_out(14) => first_stage_im_out(463),
            data_im_out(15) => first_stage_im_out(495)
        );

    ULFFT_PT16_16 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(16),
            data_re_in(1) => data_re_in(48),
            data_re_in(2) => data_re_in(80),
            data_re_in(3) => data_re_in(112),
            data_re_in(4) => data_re_in(144),
            data_re_in(5) => data_re_in(176),
            data_re_in(6) => data_re_in(208),
            data_re_in(7) => data_re_in(240),
            data_re_in(8) => data_re_in(272),
            data_re_in(9) => data_re_in(304),
            data_re_in(10) => data_re_in(336),
            data_re_in(11) => data_re_in(368),
            data_re_in(12) => data_re_in(400),
            data_re_in(13) => data_re_in(432),
            data_re_in(14) => data_re_in(464),
            data_re_in(15) => data_re_in(496),
            data_im_in(0) => data_im_in(16),
            data_im_in(1) => data_im_in(48),
            data_im_in(2) => data_im_in(80),
            data_im_in(3) => data_im_in(112),
            data_im_in(4) => data_im_in(144),
            data_im_in(5) => data_im_in(176),
            data_im_in(6) => data_im_in(208),
            data_im_in(7) => data_im_in(240),
            data_im_in(8) => data_im_in(272),
            data_im_in(9) => data_im_in(304),
            data_im_in(10) => data_im_in(336),
            data_im_in(11) => data_im_in(368),
            data_im_in(12) => data_im_in(400),
            data_im_in(13) => data_im_in(432),
            data_im_in(14) => data_im_in(464),
            data_im_in(15) => data_im_in(496),
            data_re_out(0) => first_stage_re_out(16),
            data_re_out(1) => first_stage_re_out(48),
            data_re_out(2) => first_stage_re_out(80),
            data_re_out(3) => first_stage_re_out(112),
            data_re_out(4) => first_stage_re_out(144),
            data_re_out(5) => first_stage_re_out(176),
            data_re_out(6) => first_stage_re_out(208),
            data_re_out(7) => first_stage_re_out(240),
            data_re_out(8) => first_stage_re_out(272),
            data_re_out(9) => first_stage_re_out(304),
            data_re_out(10) => first_stage_re_out(336),
            data_re_out(11) => first_stage_re_out(368),
            data_re_out(12) => first_stage_re_out(400),
            data_re_out(13) => first_stage_re_out(432),
            data_re_out(14) => first_stage_re_out(464),
            data_re_out(15) => first_stage_re_out(496),
            data_im_out(0) => first_stage_im_out(16),
            data_im_out(1) => first_stage_im_out(48),
            data_im_out(2) => first_stage_im_out(80),
            data_im_out(3) => first_stage_im_out(112),
            data_im_out(4) => first_stage_im_out(144),
            data_im_out(5) => first_stage_im_out(176),
            data_im_out(6) => first_stage_im_out(208),
            data_im_out(7) => first_stage_im_out(240),
            data_im_out(8) => first_stage_im_out(272),
            data_im_out(9) => first_stage_im_out(304),
            data_im_out(10) => first_stage_im_out(336),
            data_im_out(11) => first_stage_im_out(368),
            data_im_out(12) => first_stage_im_out(400),
            data_im_out(13) => first_stage_im_out(432),
            data_im_out(14) => first_stage_im_out(464),
            data_im_out(15) => first_stage_im_out(496)
        );

    ULFFT_PT16_17 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(17),
            data_re_in(1) => data_re_in(49),
            data_re_in(2) => data_re_in(81),
            data_re_in(3) => data_re_in(113),
            data_re_in(4) => data_re_in(145),
            data_re_in(5) => data_re_in(177),
            data_re_in(6) => data_re_in(209),
            data_re_in(7) => data_re_in(241),
            data_re_in(8) => data_re_in(273),
            data_re_in(9) => data_re_in(305),
            data_re_in(10) => data_re_in(337),
            data_re_in(11) => data_re_in(369),
            data_re_in(12) => data_re_in(401),
            data_re_in(13) => data_re_in(433),
            data_re_in(14) => data_re_in(465),
            data_re_in(15) => data_re_in(497),
            data_im_in(0) => data_im_in(17),
            data_im_in(1) => data_im_in(49),
            data_im_in(2) => data_im_in(81),
            data_im_in(3) => data_im_in(113),
            data_im_in(4) => data_im_in(145),
            data_im_in(5) => data_im_in(177),
            data_im_in(6) => data_im_in(209),
            data_im_in(7) => data_im_in(241),
            data_im_in(8) => data_im_in(273),
            data_im_in(9) => data_im_in(305),
            data_im_in(10) => data_im_in(337),
            data_im_in(11) => data_im_in(369),
            data_im_in(12) => data_im_in(401),
            data_im_in(13) => data_im_in(433),
            data_im_in(14) => data_im_in(465),
            data_im_in(15) => data_im_in(497),
            data_re_out(0) => first_stage_re_out(17),
            data_re_out(1) => first_stage_re_out(49),
            data_re_out(2) => first_stage_re_out(81),
            data_re_out(3) => first_stage_re_out(113),
            data_re_out(4) => first_stage_re_out(145),
            data_re_out(5) => first_stage_re_out(177),
            data_re_out(6) => first_stage_re_out(209),
            data_re_out(7) => first_stage_re_out(241),
            data_re_out(8) => first_stage_re_out(273),
            data_re_out(9) => first_stage_re_out(305),
            data_re_out(10) => first_stage_re_out(337),
            data_re_out(11) => first_stage_re_out(369),
            data_re_out(12) => first_stage_re_out(401),
            data_re_out(13) => first_stage_re_out(433),
            data_re_out(14) => first_stage_re_out(465),
            data_re_out(15) => first_stage_re_out(497),
            data_im_out(0) => first_stage_im_out(17),
            data_im_out(1) => first_stage_im_out(49),
            data_im_out(2) => first_stage_im_out(81),
            data_im_out(3) => first_stage_im_out(113),
            data_im_out(4) => first_stage_im_out(145),
            data_im_out(5) => first_stage_im_out(177),
            data_im_out(6) => first_stage_im_out(209),
            data_im_out(7) => first_stage_im_out(241),
            data_im_out(8) => first_stage_im_out(273),
            data_im_out(9) => first_stage_im_out(305),
            data_im_out(10) => first_stage_im_out(337),
            data_im_out(11) => first_stage_im_out(369),
            data_im_out(12) => first_stage_im_out(401),
            data_im_out(13) => first_stage_im_out(433),
            data_im_out(14) => first_stage_im_out(465),
            data_im_out(15) => first_stage_im_out(497)
        );

    ULFFT_PT16_18 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(18),
            data_re_in(1) => data_re_in(50),
            data_re_in(2) => data_re_in(82),
            data_re_in(3) => data_re_in(114),
            data_re_in(4) => data_re_in(146),
            data_re_in(5) => data_re_in(178),
            data_re_in(6) => data_re_in(210),
            data_re_in(7) => data_re_in(242),
            data_re_in(8) => data_re_in(274),
            data_re_in(9) => data_re_in(306),
            data_re_in(10) => data_re_in(338),
            data_re_in(11) => data_re_in(370),
            data_re_in(12) => data_re_in(402),
            data_re_in(13) => data_re_in(434),
            data_re_in(14) => data_re_in(466),
            data_re_in(15) => data_re_in(498),
            data_im_in(0) => data_im_in(18),
            data_im_in(1) => data_im_in(50),
            data_im_in(2) => data_im_in(82),
            data_im_in(3) => data_im_in(114),
            data_im_in(4) => data_im_in(146),
            data_im_in(5) => data_im_in(178),
            data_im_in(6) => data_im_in(210),
            data_im_in(7) => data_im_in(242),
            data_im_in(8) => data_im_in(274),
            data_im_in(9) => data_im_in(306),
            data_im_in(10) => data_im_in(338),
            data_im_in(11) => data_im_in(370),
            data_im_in(12) => data_im_in(402),
            data_im_in(13) => data_im_in(434),
            data_im_in(14) => data_im_in(466),
            data_im_in(15) => data_im_in(498),
            data_re_out(0) => first_stage_re_out(18),
            data_re_out(1) => first_stage_re_out(50),
            data_re_out(2) => first_stage_re_out(82),
            data_re_out(3) => first_stage_re_out(114),
            data_re_out(4) => first_stage_re_out(146),
            data_re_out(5) => first_stage_re_out(178),
            data_re_out(6) => first_stage_re_out(210),
            data_re_out(7) => first_stage_re_out(242),
            data_re_out(8) => first_stage_re_out(274),
            data_re_out(9) => first_stage_re_out(306),
            data_re_out(10) => first_stage_re_out(338),
            data_re_out(11) => first_stage_re_out(370),
            data_re_out(12) => first_stage_re_out(402),
            data_re_out(13) => first_stage_re_out(434),
            data_re_out(14) => first_stage_re_out(466),
            data_re_out(15) => first_stage_re_out(498),
            data_im_out(0) => first_stage_im_out(18),
            data_im_out(1) => first_stage_im_out(50),
            data_im_out(2) => first_stage_im_out(82),
            data_im_out(3) => first_stage_im_out(114),
            data_im_out(4) => first_stage_im_out(146),
            data_im_out(5) => first_stage_im_out(178),
            data_im_out(6) => first_stage_im_out(210),
            data_im_out(7) => first_stage_im_out(242),
            data_im_out(8) => first_stage_im_out(274),
            data_im_out(9) => first_stage_im_out(306),
            data_im_out(10) => first_stage_im_out(338),
            data_im_out(11) => first_stage_im_out(370),
            data_im_out(12) => first_stage_im_out(402),
            data_im_out(13) => first_stage_im_out(434),
            data_im_out(14) => first_stage_im_out(466),
            data_im_out(15) => first_stage_im_out(498)
        );

    ULFFT_PT16_19 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(19),
            data_re_in(1) => data_re_in(51),
            data_re_in(2) => data_re_in(83),
            data_re_in(3) => data_re_in(115),
            data_re_in(4) => data_re_in(147),
            data_re_in(5) => data_re_in(179),
            data_re_in(6) => data_re_in(211),
            data_re_in(7) => data_re_in(243),
            data_re_in(8) => data_re_in(275),
            data_re_in(9) => data_re_in(307),
            data_re_in(10) => data_re_in(339),
            data_re_in(11) => data_re_in(371),
            data_re_in(12) => data_re_in(403),
            data_re_in(13) => data_re_in(435),
            data_re_in(14) => data_re_in(467),
            data_re_in(15) => data_re_in(499),
            data_im_in(0) => data_im_in(19),
            data_im_in(1) => data_im_in(51),
            data_im_in(2) => data_im_in(83),
            data_im_in(3) => data_im_in(115),
            data_im_in(4) => data_im_in(147),
            data_im_in(5) => data_im_in(179),
            data_im_in(6) => data_im_in(211),
            data_im_in(7) => data_im_in(243),
            data_im_in(8) => data_im_in(275),
            data_im_in(9) => data_im_in(307),
            data_im_in(10) => data_im_in(339),
            data_im_in(11) => data_im_in(371),
            data_im_in(12) => data_im_in(403),
            data_im_in(13) => data_im_in(435),
            data_im_in(14) => data_im_in(467),
            data_im_in(15) => data_im_in(499),
            data_re_out(0) => first_stage_re_out(19),
            data_re_out(1) => first_stage_re_out(51),
            data_re_out(2) => first_stage_re_out(83),
            data_re_out(3) => first_stage_re_out(115),
            data_re_out(4) => first_stage_re_out(147),
            data_re_out(5) => first_stage_re_out(179),
            data_re_out(6) => first_stage_re_out(211),
            data_re_out(7) => first_stage_re_out(243),
            data_re_out(8) => first_stage_re_out(275),
            data_re_out(9) => first_stage_re_out(307),
            data_re_out(10) => first_stage_re_out(339),
            data_re_out(11) => first_stage_re_out(371),
            data_re_out(12) => first_stage_re_out(403),
            data_re_out(13) => first_stage_re_out(435),
            data_re_out(14) => first_stage_re_out(467),
            data_re_out(15) => first_stage_re_out(499),
            data_im_out(0) => first_stage_im_out(19),
            data_im_out(1) => first_stage_im_out(51),
            data_im_out(2) => first_stage_im_out(83),
            data_im_out(3) => first_stage_im_out(115),
            data_im_out(4) => first_stage_im_out(147),
            data_im_out(5) => first_stage_im_out(179),
            data_im_out(6) => first_stage_im_out(211),
            data_im_out(7) => first_stage_im_out(243),
            data_im_out(8) => first_stage_im_out(275),
            data_im_out(9) => first_stage_im_out(307),
            data_im_out(10) => first_stage_im_out(339),
            data_im_out(11) => first_stage_im_out(371),
            data_im_out(12) => first_stage_im_out(403),
            data_im_out(13) => first_stage_im_out(435),
            data_im_out(14) => first_stage_im_out(467),
            data_im_out(15) => first_stage_im_out(499)
        );

    ULFFT_PT16_20 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(20),
            data_re_in(1) => data_re_in(52),
            data_re_in(2) => data_re_in(84),
            data_re_in(3) => data_re_in(116),
            data_re_in(4) => data_re_in(148),
            data_re_in(5) => data_re_in(180),
            data_re_in(6) => data_re_in(212),
            data_re_in(7) => data_re_in(244),
            data_re_in(8) => data_re_in(276),
            data_re_in(9) => data_re_in(308),
            data_re_in(10) => data_re_in(340),
            data_re_in(11) => data_re_in(372),
            data_re_in(12) => data_re_in(404),
            data_re_in(13) => data_re_in(436),
            data_re_in(14) => data_re_in(468),
            data_re_in(15) => data_re_in(500),
            data_im_in(0) => data_im_in(20),
            data_im_in(1) => data_im_in(52),
            data_im_in(2) => data_im_in(84),
            data_im_in(3) => data_im_in(116),
            data_im_in(4) => data_im_in(148),
            data_im_in(5) => data_im_in(180),
            data_im_in(6) => data_im_in(212),
            data_im_in(7) => data_im_in(244),
            data_im_in(8) => data_im_in(276),
            data_im_in(9) => data_im_in(308),
            data_im_in(10) => data_im_in(340),
            data_im_in(11) => data_im_in(372),
            data_im_in(12) => data_im_in(404),
            data_im_in(13) => data_im_in(436),
            data_im_in(14) => data_im_in(468),
            data_im_in(15) => data_im_in(500),
            data_re_out(0) => first_stage_re_out(20),
            data_re_out(1) => first_stage_re_out(52),
            data_re_out(2) => first_stage_re_out(84),
            data_re_out(3) => first_stage_re_out(116),
            data_re_out(4) => first_stage_re_out(148),
            data_re_out(5) => first_stage_re_out(180),
            data_re_out(6) => first_stage_re_out(212),
            data_re_out(7) => first_stage_re_out(244),
            data_re_out(8) => first_stage_re_out(276),
            data_re_out(9) => first_stage_re_out(308),
            data_re_out(10) => first_stage_re_out(340),
            data_re_out(11) => first_stage_re_out(372),
            data_re_out(12) => first_stage_re_out(404),
            data_re_out(13) => first_stage_re_out(436),
            data_re_out(14) => first_stage_re_out(468),
            data_re_out(15) => first_stage_re_out(500),
            data_im_out(0) => first_stage_im_out(20),
            data_im_out(1) => first_stage_im_out(52),
            data_im_out(2) => first_stage_im_out(84),
            data_im_out(3) => first_stage_im_out(116),
            data_im_out(4) => first_stage_im_out(148),
            data_im_out(5) => first_stage_im_out(180),
            data_im_out(6) => first_stage_im_out(212),
            data_im_out(7) => first_stage_im_out(244),
            data_im_out(8) => first_stage_im_out(276),
            data_im_out(9) => first_stage_im_out(308),
            data_im_out(10) => first_stage_im_out(340),
            data_im_out(11) => first_stage_im_out(372),
            data_im_out(12) => first_stage_im_out(404),
            data_im_out(13) => first_stage_im_out(436),
            data_im_out(14) => first_stage_im_out(468),
            data_im_out(15) => first_stage_im_out(500)
        );

    ULFFT_PT16_21 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(21),
            data_re_in(1) => data_re_in(53),
            data_re_in(2) => data_re_in(85),
            data_re_in(3) => data_re_in(117),
            data_re_in(4) => data_re_in(149),
            data_re_in(5) => data_re_in(181),
            data_re_in(6) => data_re_in(213),
            data_re_in(7) => data_re_in(245),
            data_re_in(8) => data_re_in(277),
            data_re_in(9) => data_re_in(309),
            data_re_in(10) => data_re_in(341),
            data_re_in(11) => data_re_in(373),
            data_re_in(12) => data_re_in(405),
            data_re_in(13) => data_re_in(437),
            data_re_in(14) => data_re_in(469),
            data_re_in(15) => data_re_in(501),
            data_im_in(0) => data_im_in(21),
            data_im_in(1) => data_im_in(53),
            data_im_in(2) => data_im_in(85),
            data_im_in(3) => data_im_in(117),
            data_im_in(4) => data_im_in(149),
            data_im_in(5) => data_im_in(181),
            data_im_in(6) => data_im_in(213),
            data_im_in(7) => data_im_in(245),
            data_im_in(8) => data_im_in(277),
            data_im_in(9) => data_im_in(309),
            data_im_in(10) => data_im_in(341),
            data_im_in(11) => data_im_in(373),
            data_im_in(12) => data_im_in(405),
            data_im_in(13) => data_im_in(437),
            data_im_in(14) => data_im_in(469),
            data_im_in(15) => data_im_in(501),
            data_re_out(0) => first_stage_re_out(21),
            data_re_out(1) => first_stage_re_out(53),
            data_re_out(2) => first_stage_re_out(85),
            data_re_out(3) => first_stage_re_out(117),
            data_re_out(4) => first_stage_re_out(149),
            data_re_out(5) => first_stage_re_out(181),
            data_re_out(6) => first_stage_re_out(213),
            data_re_out(7) => first_stage_re_out(245),
            data_re_out(8) => first_stage_re_out(277),
            data_re_out(9) => first_stage_re_out(309),
            data_re_out(10) => first_stage_re_out(341),
            data_re_out(11) => first_stage_re_out(373),
            data_re_out(12) => first_stage_re_out(405),
            data_re_out(13) => first_stage_re_out(437),
            data_re_out(14) => first_stage_re_out(469),
            data_re_out(15) => first_stage_re_out(501),
            data_im_out(0) => first_stage_im_out(21),
            data_im_out(1) => first_stage_im_out(53),
            data_im_out(2) => first_stage_im_out(85),
            data_im_out(3) => first_stage_im_out(117),
            data_im_out(4) => first_stage_im_out(149),
            data_im_out(5) => first_stage_im_out(181),
            data_im_out(6) => first_stage_im_out(213),
            data_im_out(7) => first_stage_im_out(245),
            data_im_out(8) => first_stage_im_out(277),
            data_im_out(9) => first_stage_im_out(309),
            data_im_out(10) => first_stage_im_out(341),
            data_im_out(11) => first_stage_im_out(373),
            data_im_out(12) => first_stage_im_out(405),
            data_im_out(13) => first_stage_im_out(437),
            data_im_out(14) => first_stage_im_out(469),
            data_im_out(15) => first_stage_im_out(501)
        );

    ULFFT_PT16_22 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(22),
            data_re_in(1) => data_re_in(54),
            data_re_in(2) => data_re_in(86),
            data_re_in(3) => data_re_in(118),
            data_re_in(4) => data_re_in(150),
            data_re_in(5) => data_re_in(182),
            data_re_in(6) => data_re_in(214),
            data_re_in(7) => data_re_in(246),
            data_re_in(8) => data_re_in(278),
            data_re_in(9) => data_re_in(310),
            data_re_in(10) => data_re_in(342),
            data_re_in(11) => data_re_in(374),
            data_re_in(12) => data_re_in(406),
            data_re_in(13) => data_re_in(438),
            data_re_in(14) => data_re_in(470),
            data_re_in(15) => data_re_in(502),
            data_im_in(0) => data_im_in(22),
            data_im_in(1) => data_im_in(54),
            data_im_in(2) => data_im_in(86),
            data_im_in(3) => data_im_in(118),
            data_im_in(4) => data_im_in(150),
            data_im_in(5) => data_im_in(182),
            data_im_in(6) => data_im_in(214),
            data_im_in(7) => data_im_in(246),
            data_im_in(8) => data_im_in(278),
            data_im_in(9) => data_im_in(310),
            data_im_in(10) => data_im_in(342),
            data_im_in(11) => data_im_in(374),
            data_im_in(12) => data_im_in(406),
            data_im_in(13) => data_im_in(438),
            data_im_in(14) => data_im_in(470),
            data_im_in(15) => data_im_in(502),
            data_re_out(0) => first_stage_re_out(22),
            data_re_out(1) => first_stage_re_out(54),
            data_re_out(2) => first_stage_re_out(86),
            data_re_out(3) => first_stage_re_out(118),
            data_re_out(4) => first_stage_re_out(150),
            data_re_out(5) => first_stage_re_out(182),
            data_re_out(6) => first_stage_re_out(214),
            data_re_out(7) => first_stage_re_out(246),
            data_re_out(8) => first_stage_re_out(278),
            data_re_out(9) => first_stage_re_out(310),
            data_re_out(10) => first_stage_re_out(342),
            data_re_out(11) => first_stage_re_out(374),
            data_re_out(12) => first_stage_re_out(406),
            data_re_out(13) => first_stage_re_out(438),
            data_re_out(14) => first_stage_re_out(470),
            data_re_out(15) => first_stage_re_out(502),
            data_im_out(0) => first_stage_im_out(22),
            data_im_out(1) => first_stage_im_out(54),
            data_im_out(2) => first_stage_im_out(86),
            data_im_out(3) => first_stage_im_out(118),
            data_im_out(4) => first_stage_im_out(150),
            data_im_out(5) => first_stage_im_out(182),
            data_im_out(6) => first_stage_im_out(214),
            data_im_out(7) => first_stage_im_out(246),
            data_im_out(8) => first_stage_im_out(278),
            data_im_out(9) => first_stage_im_out(310),
            data_im_out(10) => first_stage_im_out(342),
            data_im_out(11) => first_stage_im_out(374),
            data_im_out(12) => first_stage_im_out(406),
            data_im_out(13) => first_stage_im_out(438),
            data_im_out(14) => first_stage_im_out(470),
            data_im_out(15) => first_stage_im_out(502)
        );

    ULFFT_PT16_23 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(23),
            data_re_in(1) => data_re_in(55),
            data_re_in(2) => data_re_in(87),
            data_re_in(3) => data_re_in(119),
            data_re_in(4) => data_re_in(151),
            data_re_in(5) => data_re_in(183),
            data_re_in(6) => data_re_in(215),
            data_re_in(7) => data_re_in(247),
            data_re_in(8) => data_re_in(279),
            data_re_in(9) => data_re_in(311),
            data_re_in(10) => data_re_in(343),
            data_re_in(11) => data_re_in(375),
            data_re_in(12) => data_re_in(407),
            data_re_in(13) => data_re_in(439),
            data_re_in(14) => data_re_in(471),
            data_re_in(15) => data_re_in(503),
            data_im_in(0) => data_im_in(23),
            data_im_in(1) => data_im_in(55),
            data_im_in(2) => data_im_in(87),
            data_im_in(3) => data_im_in(119),
            data_im_in(4) => data_im_in(151),
            data_im_in(5) => data_im_in(183),
            data_im_in(6) => data_im_in(215),
            data_im_in(7) => data_im_in(247),
            data_im_in(8) => data_im_in(279),
            data_im_in(9) => data_im_in(311),
            data_im_in(10) => data_im_in(343),
            data_im_in(11) => data_im_in(375),
            data_im_in(12) => data_im_in(407),
            data_im_in(13) => data_im_in(439),
            data_im_in(14) => data_im_in(471),
            data_im_in(15) => data_im_in(503),
            data_re_out(0) => first_stage_re_out(23),
            data_re_out(1) => first_stage_re_out(55),
            data_re_out(2) => first_stage_re_out(87),
            data_re_out(3) => first_stage_re_out(119),
            data_re_out(4) => first_stage_re_out(151),
            data_re_out(5) => first_stage_re_out(183),
            data_re_out(6) => first_stage_re_out(215),
            data_re_out(7) => first_stage_re_out(247),
            data_re_out(8) => first_stage_re_out(279),
            data_re_out(9) => first_stage_re_out(311),
            data_re_out(10) => first_stage_re_out(343),
            data_re_out(11) => first_stage_re_out(375),
            data_re_out(12) => first_stage_re_out(407),
            data_re_out(13) => first_stage_re_out(439),
            data_re_out(14) => first_stage_re_out(471),
            data_re_out(15) => first_stage_re_out(503),
            data_im_out(0) => first_stage_im_out(23),
            data_im_out(1) => first_stage_im_out(55),
            data_im_out(2) => first_stage_im_out(87),
            data_im_out(3) => first_stage_im_out(119),
            data_im_out(4) => first_stage_im_out(151),
            data_im_out(5) => first_stage_im_out(183),
            data_im_out(6) => first_stage_im_out(215),
            data_im_out(7) => first_stage_im_out(247),
            data_im_out(8) => first_stage_im_out(279),
            data_im_out(9) => first_stage_im_out(311),
            data_im_out(10) => first_stage_im_out(343),
            data_im_out(11) => first_stage_im_out(375),
            data_im_out(12) => first_stage_im_out(407),
            data_im_out(13) => first_stage_im_out(439),
            data_im_out(14) => first_stage_im_out(471),
            data_im_out(15) => first_stage_im_out(503)
        );

    ULFFT_PT16_24 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(24),
            data_re_in(1) => data_re_in(56),
            data_re_in(2) => data_re_in(88),
            data_re_in(3) => data_re_in(120),
            data_re_in(4) => data_re_in(152),
            data_re_in(5) => data_re_in(184),
            data_re_in(6) => data_re_in(216),
            data_re_in(7) => data_re_in(248),
            data_re_in(8) => data_re_in(280),
            data_re_in(9) => data_re_in(312),
            data_re_in(10) => data_re_in(344),
            data_re_in(11) => data_re_in(376),
            data_re_in(12) => data_re_in(408),
            data_re_in(13) => data_re_in(440),
            data_re_in(14) => data_re_in(472),
            data_re_in(15) => data_re_in(504),
            data_im_in(0) => data_im_in(24),
            data_im_in(1) => data_im_in(56),
            data_im_in(2) => data_im_in(88),
            data_im_in(3) => data_im_in(120),
            data_im_in(4) => data_im_in(152),
            data_im_in(5) => data_im_in(184),
            data_im_in(6) => data_im_in(216),
            data_im_in(7) => data_im_in(248),
            data_im_in(8) => data_im_in(280),
            data_im_in(9) => data_im_in(312),
            data_im_in(10) => data_im_in(344),
            data_im_in(11) => data_im_in(376),
            data_im_in(12) => data_im_in(408),
            data_im_in(13) => data_im_in(440),
            data_im_in(14) => data_im_in(472),
            data_im_in(15) => data_im_in(504),
            data_re_out(0) => first_stage_re_out(24),
            data_re_out(1) => first_stage_re_out(56),
            data_re_out(2) => first_stage_re_out(88),
            data_re_out(3) => first_stage_re_out(120),
            data_re_out(4) => first_stage_re_out(152),
            data_re_out(5) => first_stage_re_out(184),
            data_re_out(6) => first_stage_re_out(216),
            data_re_out(7) => first_stage_re_out(248),
            data_re_out(8) => first_stage_re_out(280),
            data_re_out(9) => first_stage_re_out(312),
            data_re_out(10) => first_stage_re_out(344),
            data_re_out(11) => first_stage_re_out(376),
            data_re_out(12) => first_stage_re_out(408),
            data_re_out(13) => first_stage_re_out(440),
            data_re_out(14) => first_stage_re_out(472),
            data_re_out(15) => first_stage_re_out(504),
            data_im_out(0) => first_stage_im_out(24),
            data_im_out(1) => first_stage_im_out(56),
            data_im_out(2) => first_stage_im_out(88),
            data_im_out(3) => first_stage_im_out(120),
            data_im_out(4) => first_stage_im_out(152),
            data_im_out(5) => first_stage_im_out(184),
            data_im_out(6) => first_stage_im_out(216),
            data_im_out(7) => first_stage_im_out(248),
            data_im_out(8) => first_stage_im_out(280),
            data_im_out(9) => first_stage_im_out(312),
            data_im_out(10) => first_stage_im_out(344),
            data_im_out(11) => first_stage_im_out(376),
            data_im_out(12) => first_stage_im_out(408),
            data_im_out(13) => first_stage_im_out(440),
            data_im_out(14) => first_stage_im_out(472),
            data_im_out(15) => first_stage_im_out(504)
        );

    ULFFT_PT16_25 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(25),
            data_re_in(1) => data_re_in(57),
            data_re_in(2) => data_re_in(89),
            data_re_in(3) => data_re_in(121),
            data_re_in(4) => data_re_in(153),
            data_re_in(5) => data_re_in(185),
            data_re_in(6) => data_re_in(217),
            data_re_in(7) => data_re_in(249),
            data_re_in(8) => data_re_in(281),
            data_re_in(9) => data_re_in(313),
            data_re_in(10) => data_re_in(345),
            data_re_in(11) => data_re_in(377),
            data_re_in(12) => data_re_in(409),
            data_re_in(13) => data_re_in(441),
            data_re_in(14) => data_re_in(473),
            data_re_in(15) => data_re_in(505),
            data_im_in(0) => data_im_in(25),
            data_im_in(1) => data_im_in(57),
            data_im_in(2) => data_im_in(89),
            data_im_in(3) => data_im_in(121),
            data_im_in(4) => data_im_in(153),
            data_im_in(5) => data_im_in(185),
            data_im_in(6) => data_im_in(217),
            data_im_in(7) => data_im_in(249),
            data_im_in(8) => data_im_in(281),
            data_im_in(9) => data_im_in(313),
            data_im_in(10) => data_im_in(345),
            data_im_in(11) => data_im_in(377),
            data_im_in(12) => data_im_in(409),
            data_im_in(13) => data_im_in(441),
            data_im_in(14) => data_im_in(473),
            data_im_in(15) => data_im_in(505),
            data_re_out(0) => first_stage_re_out(25),
            data_re_out(1) => first_stage_re_out(57),
            data_re_out(2) => first_stage_re_out(89),
            data_re_out(3) => first_stage_re_out(121),
            data_re_out(4) => first_stage_re_out(153),
            data_re_out(5) => first_stage_re_out(185),
            data_re_out(6) => first_stage_re_out(217),
            data_re_out(7) => first_stage_re_out(249),
            data_re_out(8) => first_stage_re_out(281),
            data_re_out(9) => first_stage_re_out(313),
            data_re_out(10) => first_stage_re_out(345),
            data_re_out(11) => first_stage_re_out(377),
            data_re_out(12) => first_stage_re_out(409),
            data_re_out(13) => first_stage_re_out(441),
            data_re_out(14) => first_stage_re_out(473),
            data_re_out(15) => first_stage_re_out(505),
            data_im_out(0) => first_stage_im_out(25),
            data_im_out(1) => first_stage_im_out(57),
            data_im_out(2) => first_stage_im_out(89),
            data_im_out(3) => first_stage_im_out(121),
            data_im_out(4) => first_stage_im_out(153),
            data_im_out(5) => first_stage_im_out(185),
            data_im_out(6) => first_stage_im_out(217),
            data_im_out(7) => first_stage_im_out(249),
            data_im_out(8) => first_stage_im_out(281),
            data_im_out(9) => first_stage_im_out(313),
            data_im_out(10) => first_stage_im_out(345),
            data_im_out(11) => first_stage_im_out(377),
            data_im_out(12) => first_stage_im_out(409),
            data_im_out(13) => first_stage_im_out(441),
            data_im_out(14) => first_stage_im_out(473),
            data_im_out(15) => first_stage_im_out(505)
        );

    ULFFT_PT16_26 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(26),
            data_re_in(1) => data_re_in(58),
            data_re_in(2) => data_re_in(90),
            data_re_in(3) => data_re_in(122),
            data_re_in(4) => data_re_in(154),
            data_re_in(5) => data_re_in(186),
            data_re_in(6) => data_re_in(218),
            data_re_in(7) => data_re_in(250),
            data_re_in(8) => data_re_in(282),
            data_re_in(9) => data_re_in(314),
            data_re_in(10) => data_re_in(346),
            data_re_in(11) => data_re_in(378),
            data_re_in(12) => data_re_in(410),
            data_re_in(13) => data_re_in(442),
            data_re_in(14) => data_re_in(474),
            data_re_in(15) => data_re_in(506),
            data_im_in(0) => data_im_in(26),
            data_im_in(1) => data_im_in(58),
            data_im_in(2) => data_im_in(90),
            data_im_in(3) => data_im_in(122),
            data_im_in(4) => data_im_in(154),
            data_im_in(5) => data_im_in(186),
            data_im_in(6) => data_im_in(218),
            data_im_in(7) => data_im_in(250),
            data_im_in(8) => data_im_in(282),
            data_im_in(9) => data_im_in(314),
            data_im_in(10) => data_im_in(346),
            data_im_in(11) => data_im_in(378),
            data_im_in(12) => data_im_in(410),
            data_im_in(13) => data_im_in(442),
            data_im_in(14) => data_im_in(474),
            data_im_in(15) => data_im_in(506),
            data_re_out(0) => first_stage_re_out(26),
            data_re_out(1) => first_stage_re_out(58),
            data_re_out(2) => first_stage_re_out(90),
            data_re_out(3) => first_stage_re_out(122),
            data_re_out(4) => first_stage_re_out(154),
            data_re_out(5) => first_stage_re_out(186),
            data_re_out(6) => first_stage_re_out(218),
            data_re_out(7) => first_stage_re_out(250),
            data_re_out(8) => first_stage_re_out(282),
            data_re_out(9) => first_stage_re_out(314),
            data_re_out(10) => first_stage_re_out(346),
            data_re_out(11) => first_stage_re_out(378),
            data_re_out(12) => first_stage_re_out(410),
            data_re_out(13) => first_stage_re_out(442),
            data_re_out(14) => first_stage_re_out(474),
            data_re_out(15) => first_stage_re_out(506),
            data_im_out(0) => first_stage_im_out(26),
            data_im_out(1) => first_stage_im_out(58),
            data_im_out(2) => first_stage_im_out(90),
            data_im_out(3) => first_stage_im_out(122),
            data_im_out(4) => first_stage_im_out(154),
            data_im_out(5) => first_stage_im_out(186),
            data_im_out(6) => first_stage_im_out(218),
            data_im_out(7) => first_stage_im_out(250),
            data_im_out(8) => first_stage_im_out(282),
            data_im_out(9) => first_stage_im_out(314),
            data_im_out(10) => first_stage_im_out(346),
            data_im_out(11) => first_stage_im_out(378),
            data_im_out(12) => first_stage_im_out(410),
            data_im_out(13) => first_stage_im_out(442),
            data_im_out(14) => first_stage_im_out(474),
            data_im_out(15) => first_stage_im_out(506)
        );

    ULFFT_PT16_27 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(27),
            data_re_in(1) => data_re_in(59),
            data_re_in(2) => data_re_in(91),
            data_re_in(3) => data_re_in(123),
            data_re_in(4) => data_re_in(155),
            data_re_in(5) => data_re_in(187),
            data_re_in(6) => data_re_in(219),
            data_re_in(7) => data_re_in(251),
            data_re_in(8) => data_re_in(283),
            data_re_in(9) => data_re_in(315),
            data_re_in(10) => data_re_in(347),
            data_re_in(11) => data_re_in(379),
            data_re_in(12) => data_re_in(411),
            data_re_in(13) => data_re_in(443),
            data_re_in(14) => data_re_in(475),
            data_re_in(15) => data_re_in(507),
            data_im_in(0) => data_im_in(27),
            data_im_in(1) => data_im_in(59),
            data_im_in(2) => data_im_in(91),
            data_im_in(3) => data_im_in(123),
            data_im_in(4) => data_im_in(155),
            data_im_in(5) => data_im_in(187),
            data_im_in(6) => data_im_in(219),
            data_im_in(7) => data_im_in(251),
            data_im_in(8) => data_im_in(283),
            data_im_in(9) => data_im_in(315),
            data_im_in(10) => data_im_in(347),
            data_im_in(11) => data_im_in(379),
            data_im_in(12) => data_im_in(411),
            data_im_in(13) => data_im_in(443),
            data_im_in(14) => data_im_in(475),
            data_im_in(15) => data_im_in(507),
            data_re_out(0) => first_stage_re_out(27),
            data_re_out(1) => first_stage_re_out(59),
            data_re_out(2) => first_stage_re_out(91),
            data_re_out(3) => first_stage_re_out(123),
            data_re_out(4) => first_stage_re_out(155),
            data_re_out(5) => first_stage_re_out(187),
            data_re_out(6) => first_stage_re_out(219),
            data_re_out(7) => first_stage_re_out(251),
            data_re_out(8) => first_stage_re_out(283),
            data_re_out(9) => first_stage_re_out(315),
            data_re_out(10) => first_stage_re_out(347),
            data_re_out(11) => first_stage_re_out(379),
            data_re_out(12) => first_stage_re_out(411),
            data_re_out(13) => first_stage_re_out(443),
            data_re_out(14) => first_stage_re_out(475),
            data_re_out(15) => first_stage_re_out(507),
            data_im_out(0) => first_stage_im_out(27),
            data_im_out(1) => first_stage_im_out(59),
            data_im_out(2) => first_stage_im_out(91),
            data_im_out(3) => first_stage_im_out(123),
            data_im_out(4) => first_stage_im_out(155),
            data_im_out(5) => first_stage_im_out(187),
            data_im_out(6) => first_stage_im_out(219),
            data_im_out(7) => first_stage_im_out(251),
            data_im_out(8) => first_stage_im_out(283),
            data_im_out(9) => first_stage_im_out(315),
            data_im_out(10) => first_stage_im_out(347),
            data_im_out(11) => first_stage_im_out(379),
            data_im_out(12) => first_stage_im_out(411),
            data_im_out(13) => first_stage_im_out(443),
            data_im_out(14) => first_stage_im_out(475),
            data_im_out(15) => first_stage_im_out(507)
        );

    ULFFT_PT16_28 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(28),
            data_re_in(1) => data_re_in(60),
            data_re_in(2) => data_re_in(92),
            data_re_in(3) => data_re_in(124),
            data_re_in(4) => data_re_in(156),
            data_re_in(5) => data_re_in(188),
            data_re_in(6) => data_re_in(220),
            data_re_in(7) => data_re_in(252),
            data_re_in(8) => data_re_in(284),
            data_re_in(9) => data_re_in(316),
            data_re_in(10) => data_re_in(348),
            data_re_in(11) => data_re_in(380),
            data_re_in(12) => data_re_in(412),
            data_re_in(13) => data_re_in(444),
            data_re_in(14) => data_re_in(476),
            data_re_in(15) => data_re_in(508),
            data_im_in(0) => data_im_in(28),
            data_im_in(1) => data_im_in(60),
            data_im_in(2) => data_im_in(92),
            data_im_in(3) => data_im_in(124),
            data_im_in(4) => data_im_in(156),
            data_im_in(5) => data_im_in(188),
            data_im_in(6) => data_im_in(220),
            data_im_in(7) => data_im_in(252),
            data_im_in(8) => data_im_in(284),
            data_im_in(9) => data_im_in(316),
            data_im_in(10) => data_im_in(348),
            data_im_in(11) => data_im_in(380),
            data_im_in(12) => data_im_in(412),
            data_im_in(13) => data_im_in(444),
            data_im_in(14) => data_im_in(476),
            data_im_in(15) => data_im_in(508),
            data_re_out(0) => first_stage_re_out(28),
            data_re_out(1) => first_stage_re_out(60),
            data_re_out(2) => first_stage_re_out(92),
            data_re_out(3) => first_stage_re_out(124),
            data_re_out(4) => first_stage_re_out(156),
            data_re_out(5) => first_stage_re_out(188),
            data_re_out(6) => first_stage_re_out(220),
            data_re_out(7) => first_stage_re_out(252),
            data_re_out(8) => first_stage_re_out(284),
            data_re_out(9) => first_stage_re_out(316),
            data_re_out(10) => first_stage_re_out(348),
            data_re_out(11) => first_stage_re_out(380),
            data_re_out(12) => first_stage_re_out(412),
            data_re_out(13) => first_stage_re_out(444),
            data_re_out(14) => first_stage_re_out(476),
            data_re_out(15) => first_stage_re_out(508),
            data_im_out(0) => first_stage_im_out(28),
            data_im_out(1) => first_stage_im_out(60),
            data_im_out(2) => first_stage_im_out(92),
            data_im_out(3) => first_stage_im_out(124),
            data_im_out(4) => first_stage_im_out(156),
            data_im_out(5) => first_stage_im_out(188),
            data_im_out(6) => first_stage_im_out(220),
            data_im_out(7) => first_stage_im_out(252),
            data_im_out(8) => first_stage_im_out(284),
            data_im_out(9) => first_stage_im_out(316),
            data_im_out(10) => first_stage_im_out(348),
            data_im_out(11) => first_stage_im_out(380),
            data_im_out(12) => first_stage_im_out(412),
            data_im_out(13) => first_stage_im_out(444),
            data_im_out(14) => first_stage_im_out(476),
            data_im_out(15) => first_stage_im_out(508)
        );

    ULFFT_PT16_29 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(29),
            data_re_in(1) => data_re_in(61),
            data_re_in(2) => data_re_in(93),
            data_re_in(3) => data_re_in(125),
            data_re_in(4) => data_re_in(157),
            data_re_in(5) => data_re_in(189),
            data_re_in(6) => data_re_in(221),
            data_re_in(7) => data_re_in(253),
            data_re_in(8) => data_re_in(285),
            data_re_in(9) => data_re_in(317),
            data_re_in(10) => data_re_in(349),
            data_re_in(11) => data_re_in(381),
            data_re_in(12) => data_re_in(413),
            data_re_in(13) => data_re_in(445),
            data_re_in(14) => data_re_in(477),
            data_re_in(15) => data_re_in(509),
            data_im_in(0) => data_im_in(29),
            data_im_in(1) => data_im_in(61),
            data_im_in(2) => data_im_in(93),
            data_im_in(3) => data_im_in(125),
            data_im_in(4) => data_im_in(157),
            data_im_in(5) => data_im_in(189),
            data_im_in(6) => data_im_in(221),
            data_im_in(7) => data_im_in(253),
            data_im_in(8) => data_im_in(285),
            data_im_in(9) => data_im_in(317),
            data_im_in(10) => data_im_in(349),
            data_im_in(11) => data_im_in(381),
            data_im_in(12) => data_im_in(413),
            data_im_in(13) => data_im_in(445),
            data_im_in(14) => data_im_in(477),
            data_im_in(15) => data_im_in(509),
            data_re_out(0) => first_stage_re_out(29),
            data_re_out(1) => first_stage_re_out(61),
            data_re_out(2) => first_stage_re_out(93),
            data_re_out(3) => first_stage_re_out(125),
            data_re_out(4) => first_stage_re_out(157),
            data_re_out(5) => first_stage_re_out(189),
            data_re_out(6) => first_stage_re_out(221),
            data_re_out(7) => first_stage_re_out(253),
            data_re_out(8) => first_stage_re_out(285),
            data_re_out(9) => first_stage_re_out(317),
            data_re_out(10) => first_stage_re_out(349),
            data_re_out(11) => first_stage_re_out(381),
            data_re_out(12) => first_stage_re_out(413),
            data_re_out(13) => first_stage_re_out(445),
            data_re_out(14) => first_stage_re_out(477),
            data_re_out(15) => first_stage_re_out(509),
            data_im_out(0) => first_stage_im_out(29),
            data_im_out(1) => first_stage_im_out(61),
            data_im_out(2) => first_stage_im_out(93),
            data_im_out(3) => first_stage_im_out(125),
            data_im_out(4) => first_stage_im_out(157),
            data_im_out(5) => first_stage_im_out(189),
            data_im_out(6) => first_stage_im_out(221),
            data_im_out(7) => first_stage_im_out(253),
            data_im_out(8) => first_stage_im_out(285),
            data_im_out(9) => first_stage_im_out(317),
            data_im_out(10) => first_stage_im_out(349),
            data_im_out(11) => first_stage_im_out(381),
            data_im_out(12) => first_stage_im_out(413),
            data_im_out(13) => first_stage_im_out(445),
            data_im_out(14) => first_stage_im_out(477),
            data_im_out(15) => first_stage_im_out(509)
        );

    ULFFT_PT16_30 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(30),
            data_re_in(1) => data_re_in(62),
            data_re_in(2) => data_re_in(94),
            data_re_in(3) => data_re_in(126),
            data_re_in(4) => data_re_in(158),
            data_re_in(5) => data_re_in(190),
            data_re_in(6) => data_re_in(222),
            data_re_in(7) => data_re_in(254),
            data_re_in(8) => data_re_in(286),
            data_re_in(9) => data_re_in(318),
            data_re_in(10) => data_re_in(350),
            data_re_in(11) => data_re_in(382),
            data_re_in(12) => data_re_in(414),
            data_re_in(13) => data_re_in(446),
            data_re_in(14) => data_re_in(478),
            data_re_in(15) => data_re_in(510),
            data_im_in(0) => data_im_in(30),
            data_im_in(1) => data_im_in(62),
            data_im_in(2) => data_im_in(94),
            data_im_in(3) => data_im_in(126),
            data_im_in(4) => data_im_in(158),
            data_im_in(5) => data_im_in(190),
            data_im_in(6) => data_im_in(222),
            data_im_in(7) => data_im_in(254),
            data_im_in(8) => data_im_in(286),
            data_im_in(9) => data_im_in(318),
            data_im_in(10) => data_im_in(350),
            data_im_in(11) => data_im_in(382),
            data_im_in(12) => data_im_in(414),
            data_im_in(13) => data_im_in(446),
            data_im_in(14) => data_im_in(478),
            data_im_in(15) => data_im_in(510),
            data_re_out(0) => first_stage_re_out(30),
            data_re_out(1) => first_stage_re_out(62),
            data_re_out(2) => first_stage_re_out(94),
            data_re_out(3) => first_stage_re_out(126),
            data_re_out(4) => first_stage_re_out(158),
            data_re_out(5) => first_stage_re_out(190),
            data_re_out(6) => first_stage_re_out(222),
            data_re_out(7) => first_stage_re_out(254),
            data_re_out(8) => first_stage_re_out(286),
            data_re_out(9) => first_stage_re_out(318),
            data_re_out(10) => first_stage_re_out(350),
            data_re_out(11) => first_stage_re_out(382),
            data_re_out(12) => first_stage_re_out(414),
            data_re_out(13) => first_stage_re_out(446),
            data_re_out(14) => first_stage_re_out(478),
            data_re_out(15) => first_stage_re_out(510),
            data_im_out(0) => first_stage_im_out(30),
            data_im_out(1) => first_stage_im_out(62),
            data_im_out(2) => first_stage_im_out(94),
            data_im_out(3) => first_stage_im_out(126),
            data_im_out(4) => first_stage_im_out(158),
            data_im_out(5) => first_stage_im_out(190),
            data_im_out(6) => first_stage_im_out(222),
            data_im_out(7) => first_stage_im_out(254),
            data_im_out(8) => first_stage_im_out(286),
            data_im_out(9) => first_stage_im_out(318),
            data_im_out(10) => first_stage_im_out(350),
            data_im_out(11) => first_stage_im_out(382),
            data_im_out(12) => first_stage_im_out(414),
            data_im_out(13) => first_stage_im_out(446),
            data_im_out(14) => first_stage_im_out(478),
            data_im_out(15) => first_stage_im_out(510)
        );

    ULFFT_PT16_31 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(31),
            data_re_in(1) => data_re_in(63),
            data_re_in(2) => data_re_in(95),
            data_re_in(3) => data_re_in(127),
            data_re_in(4) => data_re_in(159),
            data_re_in(5) => data_re_in(191),
            data_re_in(6) => data_re_in(223),
            data_re_in(7) => data_re_in(255),
            data_re_in(8) => data_re_in(287),
            data_re_in(9) => data_re_in(319),
            data_re_in(10) => data_re_in(351),
            data_re_in(11) => data_re_in(383),
            data_re_in(12) => data_re_in(415),
            data_re_in(13) => data_re_in(447),
            data_re_in(14) => data_re_in(479),
            data_re_in(15) => data_re_in(511),
            data_im_in(0) => data_im_in(31),
            data_im_in(1) => data_im_in(63),
            data_im_in(2) => data_im_in(95),
            data_im_in(3) => data_im_in(127),
            data_im_in(4) => data_im_in(159),
            data_im_in(5) => data_im_in(191),
            data_im_in(6) => data_im_in(223),
            data_im_in(7) => data_im_in(255),
            data_im_in(8) => data_im_in(287),
            data_im_in(9) => data_im_in(319),
            data_im_in(10) => data_im_in(351),
            data_im_in(11) => data_im_in(383),
            data_im_in(12) => data_im_in(415),
            data_im_in(13) => data_im_in(447),
            data_im_in(14) => data_im_in(479),
            data_im_in(15) => data_im_in(511),
            data_re_out(0) => first_stage_re_out(31),
            data_re_out(1) => first_stage_re_out(63),
            data_re_out(2) => first_stage_re_out(95),
            data_re_out(3) => first_stage_re_out(127),
            data_re_out(4) => first_stage_re_out(159),
            data_re_out(5) => first_stage_re_out(191),
            data_re_out(6) => first_stage_re_out(223),
            data_re_out(7) => first_stage_re_out(255),
            data_re_out(8) => first_stage_re_out(287),
            data_re_out(9) => first_stage_re_out(319),
            data_re_out(10) => first_stage_re_out(351),
            data_re_out(11) => first_stage_re_out(383),
            data_re_out(12) => first_stage_re_out(415),
            data_re_out(13) => first_stage_re_out(447),
            data_re_out(14) => first_stage_re_out(479),
            data_re_out(15) => first_stage_re_out(511),
            data_im_out(0) => first_stage_im_out(31),
            data_im_out(1) => first_stage_im_out(63),
            data_im_out(2) => first_stage_im_out(95),
            data_im_out(3) => first_stage_im_out(127),
            data_im_out(4) => first_stage_im_out(159),
            data_im_out(5) => first_stage_im_out(191),
            data_im_out(6) => first_stage_im_out(223),
            data_im_out(7) => first_stage_im_out(255),
            data_im_out(8) => first_stage_im_out(287),
            data_im_out(9) => first_stage_im_out(319),
            data_im_out(10) => first_stage_im_out(351),
            data_im_out(11) => first_stage_im_out(383),
            data_im_out(12) => first_stage_im_out(415),
            data_im_out(13) => first_stage_im_out(447),
            data_im_out(14) => first_stage_im_out(479),
            data_im_out(15) => first_stage_im_out(511)
        );


    --- right-hand-side processors
    URFFT_PT32_0 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(0),
            data_re_in(1) => mul_re_out(1),
            data_re_in(2) => mul_re_out(2),
            data_re_in(3) => mul_re_out(3),
            data_re_in(4) => mul_re_out(4),
            data_re_in(5) => mul_re_out(5),
            data_re_in(6) => mul_re_out(6),
            data_re_in(7) => mul_re_out(7),
            data_re_in(8) => mul_re_out(8),
            data_re_in(9) => mul_re_out(9),
            data_re_in(10) => mul_re_out(10),
            data_re_in(11) => mul_re_out(11),
            data_re_in(12) => mul_re_out(12),
            data_re_in(13) => mul_re_out(13),
            data_re_in(14) => mul_re_out(14),
            data_re_in(15) => mul_re_out(15),
            data_re_in(16) => mul_re_out(16),
            data_re_in(17) => mul_re_out(17),
            data_re_in(18) => mul_re_out(18),
            data_re_in(19) => mul_re_out(19),
            data_re_in(20) => mul_re_out(20),
            data_re_in(21) => mul_re_out(21),
            data_re_in(22) => mul_re_out(22),
            data_re_in(23) => mul_re_out(23),
            data_re_in(24) => mul_re_out(24),
            data_re_in(25) => mul_re_out(25),
            data_re_in(26) => mul_re_out(26),
            data_re_in(27) => mul_re_out(27),
            data_re_in(28) => mul_re_out(28),
            data_re_in(29) => mul_re_out(29),
            data_re_in(30) => mul_re_out(30),
            data_re_in(31) => mul_re_out(31),
            data_im_in(0) => mul_im_out(0),
            data_im_in(1) => mul_im_out(1),
            data_im_in(2) => mul_im_out(2),
            data_im_in(3) => mul_im_out(3),
            data_im_in(4) => mul_im_out(4),
            data_im_in(5) => mul_im_out(5),
            data_im_in(6) => mul_im_out(6),
            data_im_in(7) => mul_im_out(7),
            data_im_in(8) => mul_im_out(8),
            data_im_in(9) => mul_im_out(9),
            data_im_in(10) => mul_im_out(10),
            data_im_in(11) => mul_im_out(11),
            data_im_in(12) => mul_im_out(12),
            data_im_in(13) => mul_im_out(13),
            data_im_in(14) => mul_im_out(14),
            data_im_in(15) => mul_im_out(15),
            data_im_in(16) => mul_im_out(16),
            data_im_in(17) => mul_im_out(17),
            data_im_in(18) => mul_im_out(18),
            data_im_in(19) => mul_im_out(19),
            data_im_in(20) => mul_im_out(20),
            data_im_in(21) => mul_im_out(21),
            data_im_in(22) => mul_im_out(22),
            data_im_in(23) => mul_im_out(23),
            data_im_in(24) => mul_im_out(24),
            data_im_in(25) => mul_im_out(25),
            data_im_in(26) => mul_im_out(26),
            data_im_in(27) => mul_im_out(27),
            data_im_in(28) => mul_im_out(28),
            data_im_in(29) => mul_im_out(29),
            data_im_in(30) => mul_im_out(30),
            data_im_in(31) => mul_im_out(31),
            data_re_out(0) => data_re_out(0),
            data_re_out(1) => data_re_out(16),
            data_re_out(2) => data_re_out(32),
            data_re_out(3) => data_re_out(48),
            data_re_out(4) => data_re_out(64),
            data_re_out(5) => data_re_out(80),
            data_re_out(6) => data_re_out(96),
            data_re_out(7) => data_re_out(112),
            data_re_out(8) => data_re_out(128),
            data_re_out(9) => data_re_out(144),
            data_re_out(10) => data_re_out(160),
            data_re_out(11) => data_re_out(176),
            data_re_out(12) => data_re_out(192),
            data_re_out(13) => data_re_out(208),
            data_re_out(14) => data_re_out(224),
            data_re_out(15) => data_re_out(240),
            data_re_out(16) => data_re_out(256),
            data_re_out(17) => data_re_out(272),
            data_re_out(18) => data_re_out(288),
            data_re_out(19) => data_re_out(304),
            data_re_out(20) => data_re_out(320),
            data_re_out(21) => data_re_out(336),
            data_re_out(22) => data_re_out(352),
            data_re_out(23) => data_re_out(368),
            data_re_out(24) => data_re_out(384),
            data_re_out(25) => data_re_out(400),
            data_re_out(26) => data_re_out(416),
            data_re_out(27) => data_re_out(432),
            data_re_out(28) => data_re_out(448),
            data_re_out(29) => data_re_out(464),
            data_re_out(30) => data_re_out(480),
            data_re_out(31) => data_re_out(496),
            data_im_out(0) => data_im_out(0),
            data_im_out(1) => data_im_out(16),
            data_im_out(2) => data_im_out(32),
            data_im_out(3) => data_im_out(48),
            data_im_out(4) => data_im_out(64),
            data_im_out(5) => data_im_out(80),
            data_im_out(6) => data_im_out(96),
            data_im_out(7) => data_im_out(112),
            data_im_out(8) => data_im_out(128),
            data_im_out(9) => data_im_out(144),
            data_im_out(10) => data_im_out(160),
            data_im_out(11) => data_im_out(176),
            data_im_out(12) => data_im_out(192),
            data_im_out(13) => data_im_out(208),
            data_im_out(14) => data_im_out(224),
            data_im_out(15) => data_im_out(240),
            data_im_out(16) => data_im_out(256),
            data_im_out(17) => data_im_out(272),
            data_im_out(18) => data_im_out(288),
            data_im_out(19) => data_im_out(304),
            data_im_out(20) => data_im_out(320),
            data_im_out(21) => data_im_out(336),
            data_im_out(22) => data_im_out(352),
            data_im_out(23) => data_im_out(368),
            data_im_out(24) => data_im_out(384),
            data_im_out(25) => data_im_out(400),
            data_im_out(26) => data_im_out(416),
            data_im_out(27) => data_im_out(432),
            data_im_out(28) => data_im_out(448),
            data_im_out(29) => data_im_out(464),
            data_im_out(30) => data_im_out(480),
            data_im_out(31) => data_im_out(496)
        );           

    URFFT_PT32_1 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(32),
            data_re_in(1) => mul_re_out(33),
            data_re_in(2) => mul_re_out(34),
            data_re_in(3) => mul_re_out(35),
            data_re_in(4) => mul_re_out(36),
            data_re_in(5) => mul_re_out(37),
            data_re_in(6) => mul_re_out(38),
            data_re_in(7) => mul_re_out(39),
            data_re_in(8) => mul_re_out(40),
            data_re_in(9) => mul_re_out(41),
            data_re_in(10) => mul_re_out(42),
            data_re_in(11) => mul_re_out(43),
            data_re_in(12) => mul_re_out(44),
            data_re_in(13) => mul_re_out(45),
            data_re_in(14) => mul_re_out(46),
            data_re_in(15) => mul_re_out(47),
            data_re_in(16) => mul_re_out(48),
            data_re_in(17) => mul_re_out(49),
            data_re_in(18) => mul_re_out(50),
            data_re_in(19) => mul_re_out(51),
            data_re_in(20) => mul_re_out(52),
            data_re_in(21) => mul_re_out(53),
            data_re_in(22) => mul_re_out(54),
            data_re_in(23) => mul_re_out(55),
            data_re_in(24) => mul_re_out(56),
            data_re_in(25) => mul_re_out(57),
            data_re_in(26) => mul_re_out(58),
            data_re_in(27) => mul_re_out(59),
            data_re_in(28) => mul_re_out(60),
            data_re_in(29) => mul_re_out(61),
            data_re_in(30) => mul_re_out(62),
            data_re_in(31) => mul_re_out(63),
            data_im_in(0) => mul_im_out(32),
            data_im_in(1) => mul_im_out(33),
            data_im_in(2) => mul_im_out(34),
            data_im_in(3) => mul_im_out(35),
            data_im_in(4) => mul_im_out(36),
            data_im_in(5) => mul_im_out(37),
            data_im_in(6) => mul_im_out(38),
            data_im_in(7) => mul_im_out(39),
            data_im_in(8) => mul_im_out(40),
            data_im_in(9) => mul_im_out(41),
            data_im_in(10) => mul_im_out(42),
            data_im_in(11) => mul_im_out(43),
            data_im_in(12) => mul_im_out(44),
            data_im_in(13) => mul_im_out(45),
            data_im_in(14) => mul_im_out(46),
            data_im_in(15) => mul_im_out(47),
            data_im_in(16) => mul_im_out(48),
            data_im_in(17) => mul_im_out(49),
            data_im_in(18) => mul_im_out(50),
            data_im_in(19) => mul_im_out(51),
            data_im_in(20) => mul_im_out(52),
            data_im_in(21) => mul_im_out(53),
            data_im_in(22) => mul_im_out(54),
            data_im_in(23) => mul_im_out(55),
            data_im_in(24) => mul_im_out(56),
            data_im_in(25) => mul_im_out(57),
            data_im_in(26) => mul_im_out(58),
            data_im_in(27) => mul_im_out(59),
            data_im_in(28) => mul_im_out(60),
            data_im_in(29) => mul_im_out(61),
            data_im_in(30) => mul_im_out(62),
            data_im_in(31) => mul_im_out(63),
            data_re_out(0) => data_re_out(1),
            data_re_out(1) => data_re_out(17),
            data_re_out(2) => data_re_out(33),
            data_re_out(3) => data_re_out(49),
            data_re_out(4) => data_re_out(65),
            data_re_out(5) => data_re_out(81),
            data_re_out(6) => data_re_out(97),
            data_re_out(7) => data_re_out(113),
            data_re_out(8) => data_re_out(129),
            data_re_out(9) => data_re_out(145),
            data_re_out(10) => data_re_out(161),
            data_re_out(11) => data_re_out(177),
            data_re_out(12) => data_re_out(193),
            data_re_out(13) => data_re_out(209),
            data_re_out(14) => data_re_out(225),
            data_re_out(15) => data_re_out(241),
            data_re_out(16) => data_re_out(257),
            data_re_out(17) => data_re_out(273),
            data_re_out(18) => data_re_out(289),
            data_re_out(19) => data_re_out(305),
            data_re_out(20) => data_re_out(321),
            data_re_out(21) => data_re_out(337),
            data_re_out(22) => data_re_out(353),
            data_re_out(23) => data_re_out(369),
            data_re_out(24) => data_re_out(385),
            data_re_out(25) => data_re_out(401),
            data_re_out(26) => data_re_out(417),
            data_re_out(27) => data_re_out(433),
            data_re_out(28) => data_re_out(449),
            data_re_out(29) => data_re_out(465),
            data_re_out(30) => data_re_out(481),
            data_re_out(31) => data_re_out(497),
            data_im_out(0) => data_im_out(1),
            data_im_out(1) => data_im_out(17),
            data_im_out(2) => data_im_out(33),
            data_im_out(3) => data_im_out(49),
            data_im_out(4) => data_im_out(65),
            data_im_out(5) => data_im_out(81),
            data_im_out(6) => data_im_out(97),
            data_im_out(7) => data_im_out(113),
            data_im_out(8) => data_im_out(129),
            data_im_out(9) => data_im_out(145),
            data_im_out(10) => data_im_out(161),
            data_im_out(11) => data_im_out(177),
            data_im_out(12) => data_im_out(193),
            data_im_out(13) => data_im_out(209),
            data_im_out(14) => data_im_out(225),
            data_im_out(15) => data_im_out(241),
            data_im_out(16) => data_im_out(257),
            data_im_out(17) => data_im_out(273),
            data_im_out(18) => data_im_out(289),
            data_im_out(19) => data_im_out(305),
            data_im_out(20) => data_im_out(321),
            data_im_out(21) => data_im_out(337),
            data_im_out(22) => data_im_out(353),
            data_im_out(23) => data_im_out(369),
            data_im_out(24) => data_im_out(385),
            data_im_out(25) => data_im_out(401),
            data_im_out(26) => data_im_out(417),
            data_im_out(27) => data_im_out(433),
            data_im_out(28) => data_im_out(449),
            data_im_out(29) => data_im_out(465),
            data_im_out(30) => data_im_out(481),
            data_im_out(31) => data_im_out(497)
        );           

    URFFT_PT32_2 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(64),
            data_re_in(1) => mul_re_out(65),
            data_re_in(2) => mul_re_out(66),
            data_re_in(3) => mul_re_out(67),
            data_re_in(4) => mul_re_out(68),
            data_re_in(5) => mul_re_out(69),
            data_re_in(6) => mul_re_out(70),
            data_re_in(7) => mul_re_out(71),
            data_re_in(8) => mul_re_out(72),
            data_re_in(9) => mul_re_out(73),
            data_re_in(10) => mul_re_out(74),
            data_re_in(11) => mul_re_out(75),
            data_re_in(12) => mul_re_out(76),
            data_re_in(13) => mul_re_out(77),
            data_re_in(14) => mul_re_out(78),
            data_re_in(15) => mul_re_out(79),
            data_re_in(16) => mul_re_out(80),
            data_re_in(17) => mul_re_out(81),
            data_re_in(18) => mul_re_out(82),
            data_re_in(19) => mul_re_out(83),
            data_re_in(20) => mul_re_out(84),
            data_re_in(21) => mul_re_out(85),
            data_re_in(22) => mul_re_out(86),
            data_re_in(23) => mul_re_out(87),
            data_re_in(24) => mul_re_out(88),
            data_re_in(25) => mul_re_out(89),
            data_re_in(26) => mul_re_out(90),
            data_re_in(27) => mul_re_out(91),
            data_re_in(28) => mul_re_out(92),
            data_re_in(29) => mul_re_out(93),
            data_re_in(30) => mul_re_out(94),
            data_re_in(31) => mul_re_out(95),
            data_im_in(0) => mul_im_out(64),
            data_im_in(1) => mul_im_out(65),
            data_im_in(2) => mul_im_out(66),
            data_im_in(3) => mul_im_out(67),
            data_im_in(4) => mul_im_out(68),
            data_im_in(5) => mul_im_out(69),
            data_im_in(6) => mul_im_out(70),
            data_im_in(7) => mul_im_out(71),
            data_im_in(8) => mul_im_out(72),
            data_im_in(9) => mul_im_out(73),
            data_im_in(10) => mul_im_out(74),
            data_im_in(11) => mul_im_out(75),
            data_im_in(12) => mul_im_out(76),
            data_im_in(13) => mul_im_out(77),
            data_im_in(14) => mul_im_out(78),
            data_im_in(15) => mul_im_out(79),
            data_im_in(16) => mul_im_out(80),
            data_im_in(17) => mul_im_out(81),
            data_im_in(18) => mul_im_out(82),
            data_im_in(19) => mul_im_out(83),
            data_im_in(20) => mul_im_out(84),
            data_im_in(21) => mul_im_out(85),
            data_im_in(22) => mul_im_out(86),
            data_im_in(23) => mul_im_out(87),
            data_im_in(24) => mul_im_out(88),
            data_im_in(25) => mul_im_out(89),
            data_im_in(26) => mul_im_out(90),
            data_im_in(27) => mul_im_out(91),
            data_im_in(28) => mul_im_out(92),
            data_im_in(29) => mul_im_out(93),
            data_im_in(30) => mul_im_out(94),
            data_im_in(31) => mul_im_out(95),
            data_re_out(0) => data_re_out(2),
            data_re_out(1) => data_re_out(18),
            data_re_out(2) => data_re_out(34),
            data_re_out(3) => data_re_out(50),
            data_re_out(4) => data_re_out(66),
            data_re_out(5) => data_re_out(82),
            data_re_out(6) => data_re_out(98),
            data_re_out(7) => data_re_out(114),
            data_re_out(8) => data_re_out(130),
            data_re_out(9) => data_re_out(146),
            data_re_out(10) => data_re_out(162),
            data_re_out(11) => data_re_out(178),
            data_re_out(12) => data_re_out(194),
            data_re_out(13) => data_re_out(210),
            data_re_out(14) => data_re_out(226),
            data_re_out(15) => data_re_out(242),
            data_re_out(16) => data_re_out(258),
            data_re_out(17) => data_re_out(274),
            data_re_out(18) => data_re_out(290),
            data_re_out(19) => data_re_out(306),
            data_re_out(20) => data_re_out(322),
            data_re_out(21) => data_re_out(338),
            data_re_out(22) => data_re_out(354),
            data_re_out(23) => data_re_out(370),
            data_re_out(24) => data_re_out(386),
            data_re_out(25) => data_re_out(402),
            data_re_out(26) => data_re_out(418),
            data_re_out(27) => data_re_out(434),
            data_re_out(28) => data_re_out(450),
            data_re_out(29) => data_re_out(466),
            data_re_out(30) => data_re_out(482),
            data_re_out(31) => data_re_out(498),
            data_im_out(0) => data_im_out(2),
            data_im_out(1) => data_im_out(18),
            data_im_out(2) => data_im_out(34),
            data_im_out(3) => data_im_out(50),
            data_im_out(4) => data_im_out(66),
            data_im_out(5) => data_im_out(82),
            data_im_out(6) => data_im_out(98),
            data_im_out(7) => data_im_out(114),
            data_im_out(8) => data_im_out(130),
            data_im_out(9) => data_im_out(146),
            data_im_out(10) => data_im_out(162),
            data_im_out(11) => data_im_out(178),
            data_im_out(12) => data_im_out(194),
            data_im_out(13) => data_im_out(210),
            data_im_out(14) => data_im_out(226),
            data_im_out(15) => data_im_out(242),
            data_im_out(16) => data_im_out(258),
            data_im_out(17) => data_im_out(274),
            data_im_out(18) => data_im_out(290),
            data_im_out(19) => data_im_out(306),
            data_im_out(20) => data_im_out(322),
            data_im_out(21) => data_im_out(338),
            data_im_out(22) => data_im_out(354),
            data_im_out(23) => data_im_out(370),
            data_im_out(24) => data_im_out(386),
            data_im_out(25) => data_im_out(402),
            data_im_out(26) => data_im_out(418),
            data_im_out(27) => data_im_out(434),
            data_im_out(28) => data_im_out(450),
            data_im_out(29) => data_im_out(466),
            data_im_out(30) => data_im_out(482),
            data_im_out(31) => data_im_out(498)
        );           

    URFFT_PT32_3 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(96),
            data_re_in(1) => mul_re_out(97),
            data_re_in(2) => mul_re_out(98),
            data_re_in(3) => mul_re_out(99),
            data_re_in(4) => mul_re_out(100),
            data_re_in(5) => mul_re_out(101),
            data_re_in(6) => mul_re_out(102),
            data_re_in(7) => mul_re_out(103),
            data_re_in(8) => mul_re_out(104),
            data_re_in(9) => mul_re_out(105),
            data_re_in(10) => mul_re_out(106),
            data_re_in(11) => mul_re_out(107),
            data_re_in(12) => mul_re_out(108),
            data_re_in(13) => mul_re_out(109),
            data_re_in(14) => mul_re_out(110),
            data_re_in(15) => mul_re_out(111),
            data_re_in(16) => mul_re_out(112),
            data_re_in(17) => mul_re_out(113),
            data_re_in(18) => mul_re_out(114),
            data_re_in(19) => mul_re_out(115),
            data_re_in(20) => mul_re_out(116),
            data_re_in(21) => mul_re_out(117),
            data_re_in(22) => mul_re_out(118),
            data_re_in(23) => mul_re_out(119),
            data_re_in(24) => mul_re_out(120),
            data_re_in(25) => mul_re_out(121),
            data_re_in(26) => mul_re_out(122),
            data_re_in(27) => mul_re_out(123),
            data_re_in(28) => mul_re_out(124),
            data_re_in(29) => mul_re_out(125),
            data_re_in(30) => mul_re_out(126),
            data_re_in(31) => mul_re_out(127),
            data_im_in(0) => mul_im_out(96),
            data_im_in(1) => mul_im_out(97),
            data_im_in(2) => mul_im_out(98),
            data_im_in(3) => mul_im_out(99),
            data_im_in(4) => mul_im_out(100),
            data_im_in(5) => mul_im_out(101),
            data_im_in(6) => mul_im_out(102),
            data_im_in(7) => mul_im_out(103),
            data_im_in(8) => mul_im_out(104),
            data_im_in(9) => mul_im_out(105),
            data_im_in(10) => mul_im_out(106),
            data_im_in(11) => mul_im_out(107),
            data_im_in(12) => mul_im_out(108),
            data_im_in(13) => mul_im_out(109),
            data_im_in(14) => mul_im_out(110),
            data_im_in(15) => mul_im_out(111),
            data_im_in(16) => mul_im_out(112),
            data_im_in(17) => mul_im_out(113),
            data_im_in(18) => mul_im_out(114),
            data_im_in(19) => mul_im_out(115),
            data_im_in(20) => mul_im_out(116),
            data_im_in(21) => mul_im_out(117),
            data_im_in(22) => mul_im_out(118),
            data_im_in(23) => mul_im_out(119),
            data_im_in(24) => mul_im_out(120),
            data_im_in(25) => mul_im_out(121),
            data_im_in(26) => mul_im_out(122),
            data_im_in(27) => mul_im_out(123),
            data_im_in(28) => mul_im_out(124),
            data_im_in(29) => mul_im_out(125),
            data_im_in(30) => mul_im_out(126),
            data_im_in(31) => mul_im_out(127),
            data_re_out(0) => data_re_out(3),
            data_re_out(1) => data_re_out(19),
            data_re_out(2) => data_re_out(35),
            data_re_out(3) => data_re_out(51),
            data_re_out(4) => data_re_out(67),
            data_re_out(5) => data_re_out(83),
            data_re_out(6) => data_re_out(99),
            data_re_out(7) => data_re_out(115),
            data_re_out(8) => data_re_out(131),
            data_re_out(9) => data_re_out(147),
            data_re_out(10) => data_re_out(163),
            data_re_out(11) => data_re_out(179),
            data_re_out(12) => data_re_out(195),
            data_re_out(13) => data_re_out(211),
            data_re_out(14) => data_re_out(227),
            data_re_out(15) => data_re_out(243),
            data_re_out(16) => data_re_out(259),
            data_re_out(17) => data_re_out(275),
            data_re_out(18) => data_re_out(291),
            data_re_out(19) => data_re_out(307),
            data_re_out(20) => data_re_out(323),
            data_re_out(21) => data_re_out(339),
            data_re_out(22) => data_re_out(355),
            data_re_out(23) => data_re_out(371),
            data_re_out(24) => data_re_out(387),
            data_re_out(25) => data_re_out(403),
            data_re_out(26) => data_re_out(419),
            data_re_out(27) => data_re_out(435),
            data_re_out(28) => data_re_out(451),
            data_re_out(29) => data_re_out(467),
            data_re_out(30) => data_re_out(483),
            data_re_out(31) => data_re_out(499),
            data_im_out(0) => data_im_out(3),
            data_im_out(1) => data_im_out(19),
            data_im_out(2) => data_im_out(35),
            data_im_out(3) => data_im_out(51),
            data_im_out(4) => data_im_out(67),
            data_im_out(5) => data_im_out(83),
            data_im_out(6) => data_im_out(99),
            data_im_out(7) => data_im_out(115),
            data_im_out(8) => data_im_out(131),
            data_im_out(9) => data_im_out(147),
            data_im_out(10) => data_im_out(163),
            data_im_out(11) => data_im_out(179),
            data_im_out(12) => data_im_out(195),
            data_im_out(13) => data_im_out(211),
            data_im_out(14) => data_im_out(227),
            data_im_out(15) => data_im_out(243),
            data_im_out(16) => data_im_out(259),
            data_im_out(17) => data_im_out(275),
            data_im_out(18) => data_im_out(291),
            data_im_out(19) => data_im_out(307),
            data_im_out(20) => data_im_out(323),
            data_im_out(21) => data_im_out(339),
            data_im_out(22) => data_im_out(355),
            data_im_out(23) => data_im_out(371),
            data_im_out(24) => data_im_out(387),
            data_im_out(25) => data_im_out(403),
            data_im_out(26) => data_im_out(419),
            data_im_out(27) => data_im_out(435),
            data_im_out(28) => data_im_out(451),
            data_im_out(29) => data_im_out(467),
            data_im_out(30) => data_im_out(483),
            data_im_out(31) => data_im_out(499)
        );           

    URFFT_PT32_4 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(128),
            data_re_in(1) => mul_re_out(129),
            data_re_in(2) => mul_re_out(130),
            data_re_in(3) => mul_re_out(131),
            data_re_in(4) => mul_re_out(132),
            data_re_in(5) => mul_re_out(133),
            data_re_in(6) => mul_re_out(134),
            data_re_in(7) => mul_re_out(135),
            data_re_in(8) => mul_re_out(136),
            data_re_in(9) => mul_re_out(137),
            data_re_in(10) => mul_re_out(138),
            data_re_in(11) => mul_re_out(139),
            data_re_in(12) => mul_re_out(140),
            data_re_in(13) => mul_re_out(141),
            data_re_in(14) => mul_re_out(142),
            data_re_in(15) => mul_re_out(143),
            data_re_in(16) => mul_re_out(144),
            data_re_in(17) => mul_re_out(145),
            data_re_in(18) => mul_re_out(146),
            data_re_in(19) => mul_re_out(147),
            data_re_in(20) => mul_re_out(148),
            data_re_in(21) => mul_re_out(149),
            data_re_in(22) => mul_re_out(150),
            data_re_in(23) => mul_re_out(151),
            data_re_in(24) => mul_re_out(152),
            data_re_in(25) => mul_re_out(153),
            data_re_in(26) => mul_re_out(154),
            data_re_in(27) => mul_re_out(155),
            data_re_in(28) => mul_re_out(156),
            data_re_in(29) => mul_re_out(157),
            data_re_in(30) => mul_re_out(158),
            data_re_in(31) => mul_re_out(159),
            data_im_in(0) => mul_im_out(128),
            data_im_in(1) => mul_im_out(129),
            data_im_in(2) => mul_im_out(130),
            data_im_in(3) => mul_im_out(131),
            data_im_in(4) => mul_im_out(132),
            data_im_in(5) => mul_im_out(133),
            data_im_in(6) => mul_im_out(134),
            data_im_in(7) => mul_im_out(135),
            data_im_in(8) => mul_im_out(136),
            data_im_in(9) => mul_im_out(137),
            data_im_in(10) => mul_im_out(138),
            data_im_in(11) => mul_im_out(139),
            data_im_in(12) => mul_im_out(140),
            data_im_in(13) => mul_im_out(141),
            data_im_in(14) => mul_im_out(142),
            data_im_in(15) => mul_im_out(143),
            data_im_in(16) => mul_im_out(144),
            data_im_in(17) => mul_im_out(145),
            data_im_in(18) => mul_im_out(146),
            data_im_in(19) => mul_im_out(147),
            data_im_in(20) => mul_im_out(148),
            data_im_in(21) => mul_im_out(149),
            data_im_in(22) => mul_im_out(150),
            data_im_in(23) => mul_im_out(151),
            data_im_in(24) => mul_im_out(152),
            data_im_in(25) => mul_im_out(153),
            data_im_in(26) => mul_im_out(154),
            data_im_in(27) => mul_im_out(155),
            data_im_in(28) => mul_im_out(156),
            data_im_in(29) => mul_im_out(157),
            data_im_in(30) => mul_im_out(158),
            data_im_in(31) => mul_im_out(159),
            data_re_out(0) => data_re_out(4),
            data_re_out(1) => data_re_out(20),
            data_re_out(2) => data_re_out(36),
            data_re_out(3) => data_re_out(52),
            data_re_out(4) => data_re_out(68),
            data_re_out(5) => data_re_out(84),
            data_re_out(6) => data_re_out(100),
            data_re_out(7) => data_re_out(116),
            data_re_out(8) => data_re_out(132),
            data_re_out(9) => data_re_out(148),
            data_re_out(10) => data_re_out(164),
            data_re_out(11) => data_re_out(180),
            data_re_out(12) => data_re_out(196),
            data_re_out(13) => data_re_out(212),
            data_re_out(14) => data_re_out(228),
            data_re_out(15) => data_re_out(244),
            data_re_out(16) => data_re_out(260),
            data_re_out(17) => data_re_out(276),
            data_re_out(18) => data_re_out(292),
            data_re_out(19) => data_re_out(308),
            data_re_out(20) => data_re_out(324),
            data_re_out(21) => data_re_out(340),
            data_re_out(22) => data_re_out(356),
            data_re_out(23) => data_re_out(372),
            data_re_out(24) => data_re_out(388),
            data_re_out(25) => data_re_out(404),
            data_re_out(26) => data_re_out(420),
            data_re_out(27) => data_re_out(436),
            data_re_out(28) => data_re_out(452),
            data_re_out(29) => data_re_out(468),
            data_re_out(30) => data_re_out(484),
            data_re_out(31) => data_re_out(500),
            data_im_out(0) => data_im_out(4),
            data_im_out(1) => data_im_out(20),
            data_im_out(2) => data_im_out(36),
            data_im_out(3) => data_im_out(52),
            data_im_out(4) => data_im_out(68),
            data_im_out(5) => data_im_out(84),
            data_im_out(6) => data_im_out(100),
            data_im_out(7) => data_im_out(116),
            data_im_out(8) => data_im_out(132),
            data_im_out(9) => data_im_out(148),
            data_im_out(10) => data_im_out(164),
            data_im_out(11) => data_im_out(180),
            data_im_out(12) => data_im_out(196),
            data_im_out(13) => data_im_out(212),
            data_im_out(14) => data_im_out(228),
            data_im_out(15) => data_im_out(244),
            data_im_out(16) => data_im_out(260),
            data_im_out(17) => data_im_out(276),
            data_im_out(18) => data_im_out(292),
            data_im_out(19) => data_im_out(308),
            data_im_out(20) => data_im_out(324),
            data_im_out(21) => data_im_out(340),
            data_im_out(22) => data_im_out(356),
            data_im_out(23) => data_im_out(372),
            data_im_out(24) => data_im_out(388),
            data_im_out(25) => data_im_out(404),
            data_im_out(26) => data_im_out(420),
            data_im_out(27) => data_im_out(436),
            data_im_out(28) => data_im_out(452),
            data_im_out(29) => data_im_out(468),
            data_im_out(30) => data_im_out(484),
            data_im_out(31) => data_im_out(500)
        );           

    URFFT_PT32_5 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(160),
            data_re_in(1) => mul_re_out(161),
            data_re_in(2) => mul_re_out(162),
            data_re_in(3) => mul_re_out(163),
            data_re_in(4) => mul_re_out(164),
            data_re_in(5) => mul_re_out(165),
            data_re_in(6) => mul_re_out(166),
            data_re_in(7) => mul_re_out(167),
            data_re_in(8) => mul_re_out(168),
            data_re_in(9) => mul_re_out(169),
            data_re_in(10) => mul_re_out(170),
            data_re_in(11) => mul_re_out(171),
            data_re_in(12) => mul_re_out(172),
            data_re_in(13) => mul_re_out(173),
            data_re_in(14) => mul_re_out(174),
            data_re_in(15) => mul_re_out(175),
            data_re_in(16) => mul_re_out(176),
            data_re_in(17) => mul_re_out(177),
            data_re_in(18) => mul_re_out(178),
            data_re_in(19) => mul_re_out(179),
            data_re_in(20) => mul_re_out(180),
            data_re_in(21) => mul_re_out(181),
            data_re_in(22) => mul_re_out(182),
            data_re_in(23) => mul_re_out(183),
            data_re_in(24) => mul_re_out(184),
            data_re_in(25) => mul_re_out(185),
            data_re_in(26) => mul_re_out(186),
            data_re_in(27) => mul_re_out(187),
            data_re_in(28) => mul_re_out(188),
            data_re_in(29) => mul_re_out(189),
            data_re_in(30) => mul_re_out(190),
            data_re_in(31) => mul_re_out(191),
            data_im_in(0) => mul_im_out(160),
            data_im_in(1) => mul_im_out(161),
            data_im_in(2) => mul_im_out(162),
            data_im_in(3) => mul_im_out(163),
            data_im_in(4) => mul_im_out(164),
            data_im_in(5) => mul_im_out(165),
            data_im_in(6) => mul_im_out(166),
            data_im_in(7) => mul_im_out(167),
            data_im_in(8) => mul_im_out(168),
            data_im_in(9) => mul_im_out(169),
            data_im_in(10) => mul_im_out(170),
            data_im_in(11) => mul_im_out(171),
            data_im_in(12) => mul_im_out(172),
            data_im_in(13) => mul_im_out(173),
            data_im_in(14) => mul_im_out(174),
            data_im_in(15) => mul_im_out(175),
            data_im_in(16) => mul_im_out(176),
            data_im_in(17) => mul_im_out(177),
            data_im_in(18) => mul_im_out(178),
            data_im_in(19) => mul_im_out(179),
            data_im_in(20) => mul_im_out(180),
            data_im_in(21) => mul_im_out(181),
            data_im_in(22) => mul_im_out(182),
            data_im_in(23) => mul_im_out(183),
            data_im_in(24) => mul_im_out(184),
            data_im_in(25) => mul_im_out(185),
            data_im_in(26) => mul_im_out(186),
            data_im_in(27) => mul_im_out(187),
            data_im_in(28) => mul_im_out(188),
            data_im_in(29) => mul_im_out(189),
            data_im_in(30) => mul_im_out(190),
            data_im_in(31) => mul_im_out(191),
            data_re_out(0) => data_re_out(5),
            data_re_out(1) => data_re_out(21),
            data_re_out(2) => data_re_out(37),
            data_re_out(3) => data_re_out(53),
            data_re_out(4) => data_re_out(69),
            data_re_out(5) => data_re_out(85),
            data_re_out(6) => data_re_out(101),
            data_re_out(7) => data_re_out(117),
            data_re_out(8) => data_re_out(133),
            data_re_out(9) => data_re_out(149),
            data_re_out(10) => data_re_out(165),
            data_re_out(11) => data_re_out(181),
            data_re_out(12) => data_re_out(197),
            data_re_out(13) => data_re_out(213),
            data_re_out(14) => data_re_out(229),
            data_re_out(15) => data_re_out(245),
            data_re_out(16) => data_re_out(261),
            data_re_out(17) => data_re_out(277),
            data_re_out(18) => data_re_out(293),
            data_re_out(19) => data_re_out(309),
            data_re_out(20) => data_re_out(325),
            data_re_out(21) => data_re_out(341),
            data_re_out(22) => data_re_out(357),
            data_re_out(23) => data_re_out(373),
            data_re_out(24) => data_re_out(389),
            data_re_out(25) => data_re_out(405),
            data_re_out(26) => data_re_out(421),
            data_re_out(27) => data_re_out(437),
            data_re_out(28) => data_re_out(453),
            data_re_out(29) => data_re_out(469),
            data_re_out(30) => data_re_out(485),
            data_re_out(31) => data_re_out(501),
            data_im_out(0) => data_im_out(5),
            data_im_out(1) => data_im_out(21),
            data_im_out(2) => data_im_out(37),
            data_im_out(3) => data_im_out(53),
            data_im_out(4) => data_im_out(69),
            data_im_out(5) => data_im_out(85),
            data_im_out(6) => data_im_out(101),
            data_im_out(7) => data_im_out(117),
            data_im_out(8) => data_im_out(133),
            data_im_out(9) => data_im_out(149),
            data_im_out(10) => data_im_out(165),
            data_im_out(11) => data_im_out(181),
            data_im_out(12) => data_im_out(197),
            data_im_out(13) => data_im_out(213),
            data_im_out(14) => data_im_out(229),
            data_im_out(15) => data_im_out(245),
            data_im_out(16) => data_im_out(261),
            data_im_out(17) => data_im_out(277),
            data_im_out(18) => data_im_out(293),
            data_im_out(19) => data_im_out(309),
            data_im_out(20) => data_im_out(325),
            data_im_out(21) => data_im_out(341),
            data_im_out(22) => data_im_out(357),
            data_im_out(23) => data_im_out(373),
            data_im_out(24) => data_im_out(389),
            data_im_out(25) => data_im_out(405),
            data_im_out(26) => data_im_out(421),
            data_im_out(27) => data_im_out(437),
            data_im_out(28) => data_im_out(453),
            data_im_out(29) => data_im_out(469),
            data_im_out(30) => data_im_out(485),
            data_im_out(31) => data_im_out(501)
        );           

    URFFT_PT32_6 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(192),
            data_re_in(1) => mul_re_out(193),
            data_re_in(2) => mul_re_out(194),
            data_re_in(3) => mul_re_out(195),
            data_re_in(4) => mul_re_out(196),
            data_re_in(5) => mul_re_out(197),
            data_re_in(6) => mul_re_out(198),
            data_re_in(7) => mul_re_out(199),
            data_re_in(8) => mul_re_out(200),
            data_re_in(9) => mul_re_out(201),
            data_re_in(10) => mul_re_out(202),
            data_re_in(11) => mul_re_out(203),
            data_re_in(12) => mul_re_out(204),
            data_re_in(13) => mul_re_out(205),
            data_re_in(14) => mul_re_out(206),
            data_re_in(15) => mul_re_out(207),
            data_re_in(16) => mul_re_out(208),
            data_re_in(17) => mul_re_out(209),
            data_re_in(18) => mul_re_out(210),
            data_re_in(19) => mul_re_out(211),
            data_re_in(20) => mul_re_out(212),
            data_re_in(21) => mul_re_out(213),
            data_re_in(22) => mul_re_out(214),
            data_re_in(23) => mul_re_out(215),
            data_re_in(24) => mul_re_out(216),
            data_re_in(25) => mul_re_out(217),
            data_re_in(26) => mul_re_out(218),
            data_re_in(27) => mul_re_out(219),
            data_re_in(28) => mul_re_out(220),
            data_re_in(29) => mul_re_out(221),
            data_re_in(30) => mul_re_out(222),
            data_re_in(31) => mul_re_out(223),
            data_im_in(0) => mul_im_out(192),
            data_im_in(1) => mul_im_out(193),
            data_im_in(2) => mul_im_out(194),
            data_im_in(3) => mul_im_out(195),
            data_im_in(4) => mul_im_out(196),
            data_im_in(5) => mul_im_out(197),
            data_im_in(6) => mul_im_out(198),
            data_im_in(7) => mul_im_out(199),
            data_im_in(8) => mul_im_out(200),
            data_im_in(9) => mul_im_out(201),
            data_im_in(10) => mul_im_out(202),
            data_im_in(11) => mul_im_out(203),
            data_im_in(12) => mul_im_out(204),
            data_im_in(13) => mul_im_out(205),
            data_im_in(14) => mul_im_out(206),
            data_im_in(15) => mul_im_out(207),
            data_im_in(16) => mul_im_out(208),
            data_im_in(17) => mul_im_out(209),
            data_im_in(18) => mul_im_out(210),
            data_im_in(19) => mul_im_out(211),
            data_im_in(20) => mul_im_out(212),
            data_im_in(21) => mul_im_out(213),
            data_im_in(22) => mul_im_out(214),
            data_im_in(23) => mul_im_out(215),
            data_im_in(24) => mul_im_out(216),
            data_im_in(25) => mul_im_out(217),
            data_im_in(26) => mul_im_out(218),
            data_im_in(27) => mul_im_out(219),
            data_im_in(28) => mul_im_out(220),
            data_im_in(29) => mul_im_out(221),
            data_im_in(30) => mul_im_out(222),
            data_im_in(31) => mul_im_out(223),
            data_re_out(0) => data_re_out(6),
            data_re_out(1) => data_re_out(22),
            data_re_out(2) => data_re_out(38),
            data_re_out(3) => data_re_out(54),
            data_re_out(4) => data_re_out(70),
            data_re_out(5) => data_re_out(86),
            data_re_out(6) => data_re_out(102),
            data_re_out(7) => data_re_out(118),
            data_re_out(8) => data_re_out(134),
            data_re_out(9) => data_re_out(150),
            data_re_out(10) => data_re_out(166),
            data_re_out(11) => data_re_out(182),
            data_re_out(12) => data_re_out(198),
            data_re_out(13) => data_re_out(214),
            data_re_out(14) => data_re_out(230),
            data_re_out(15) => data_re_out(246),
            data_re_out(16) => data_re_out(262),
            data_re_out(17) => data_re_out(278),
            data_re_out(18) => data_re_out(294),
            data_re_out(19) => data_re_out(310),
            data_re_out(20) => data_re_out(326),
            data_re_out(21) => data_re_out(342),
            data_re_out(22) => data_re_out(358),
            data_re_out(23) => data_re_out(374),
            data_re_out(24) => data_re_out(390),
            data_re_out(25) => data_re_out(406),
            data_re_out(26) => data_re_out(422),
            data_re_out(27) => data_re_out(438),
            data_re_out(28) => data_re_out(454),
            data_re_out(29) => data_re_out(470),
            data_re_out(30) => data_re_out(486),
            data_re_out(31) => data_re_out(502),
            data_im_out(0) => data_im_out(6),
            data_im_out(1) => data_im_out(22),
            data_im_out(2) => data_im_out(38),
            data_im_out(3) => data_im_out(54),
            data_im_out(4) => data_im_out(70),
            data_im_out(5) => data_im_out(86),
            data_im_out(6) => data_im_out(102),
            data_im_out(7) => data_im_out(118),
            data_im_out(8) => data_im_out(134),
            data_im_out(9) => data_im_out(150),
            data_im_out(10) => data_im_out(166),
            data_im_out(11) => data_im_out(182),
            data_im_out(12) => data_im_out(198),
            data_im_out(13) => data_im_out(214),
            data_im_out(14) => data_im_out(230),
            data_im_out(15) => data_im_out(246),
            data_im_out(16) => data_im_out(262),
            data_im_out(17) => data_im_out(278),
            data_im_out(18) => data_im_out(294),
            data_im_out(19) => data_im_out(310),
            data_im_out(20) => data_im_out(326),
            data_im_out(21) => data_im_out(342),
            data_im_out(22) => data_im_out(358),
            data_im_out(23) => data_im_out(374),
            data_im_out(24) => data_im_out(390),
            data_im_out(25) => data_im_out(406),
            data_im_out(26) => data_im_out(422),
            data_im_out(27) => data_im_out(438),
            data_im_out(28) => data_im_out(454),
            data_im_out(29) => data_im_out(470),
            data_im_out(30) => data_im_out(486),
            data_im_out(31) => data_im_out(502)
        );           

    URFFT_PT32_7 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(224),
            data_re_in(1) => mul_re_out(225),
            data_re_in(2) => mul_re_out(226),
            data_re_in(3) => mul_re_out(227),
            data_re_in(4) => mul_re_out(228),
            data_re_in(5) => mul_re_out(229),
            data_re_in(6) => mul_re_out(230),
            data_re_in(7) => mul_re_out(231),
            data_re_in(8) => mul_re_out(232),
            data_re_in(9) => mul_re_out(233),
            data_re_in(10) => mul_re_out(234),
            data_re_in(11) => mul_re_out(235),
            data_re_in(12) => mul_re_out(236),
            data_re_in(13) => mul_re_out(237),
            data_re_in(14) => mul_re_out(238),
            data_re_in(15) => mul_re_out(239),
            data_re_in(16) => mul_re_out(240),
            data_re_in(17) => mul_re_out(241),
            data_re_in(18) => mul_re_out(242),
            data_re_in(19) => mul_re_out(243),
            data_re_in(20) => mul_re_out(244),
            data_re_in(21) => mul_re_out(245),
            data_re_in(22) => mul_re_out(246),
            data_re_in(23) => mul_re_out(247),
            data_re_in(24) => mul_re_out(248),
            data_re_in(25) => mul_re_out(249),
            data_re_in(26) => mul_re_out(250),
            data_re_in(27) => mul_re_out(251),
            data_re_in(28) => mul_re_out(252),
            data_re_in(29) => mul_re_out(253),
            data_re_in(30) => mul_re_out(254),
            data_re_in(31) => mul_re_out(255),
            data_im_in(0) => mul_im_out(224),
            data_im_in(1) => mul_im_out(225),
            data_im_in(2) => mul_im_out(226),
            data_im_in(3) => mul_im_out(227),
            data_im_in(4) => mul_im_out(228),
            data_im_in(5) => mul_im_out(229),
            data_im_in(6) => mul_im_out(230),
            data_im_in(7) => mul_im_out(231),
            data_im_in(8) => mul_im_out(232),
            data_im_in(9) => mul_im_out(233),
            data_im_in(10) => mul_im_out(234),
            data_im_in(11) => mul_im_out(235),
            data_im_in(12) => mul_im_out(236),
            data_im_in(13) => mul_im_out(237),
            data_im_in(14) => mul_im_out(238),
            data_im_in(15) => mul_im_out(239),
            data_im_in(16) => mul_im_out(240),
            data_im_in(17) => mul_im_out(241),
            data_im_in(18) => mul_im_out(242),
            data_im_in(19) => mul_im_out(243),
            data_im_in(20) => mul_im_out(244),
            data_im_in(21) => mul_im_out(245),
            data_im_in(22) => mul_im_out(246),
            data_im_in(23) => mul_im_out(247),
            data_im_in(24) => mul_im_out(248),
            data_im_in(25) => mul_im_out(249),
            data_im_in(26) => mul_im_out(250),
            data_im_in(27) => mul_im_out(251),
            data_im_in(28) => mul_im_out(252),
            data_im_in(29) => mul_im_out(253),
            data_im_in(30) => mul_im_out(254),
            data_im_in(31) => mul_im_out(255),
            data_re_out(0) => data_re_out(7),
            data_re_out(1) => data_re_out(23),
            data_re_out(2) => data_re_out(39),
            data_re_out(3) => data_re_out(55),
            data_re_out(4) => data_re_out(71),
            data_re_out(5) => data_re_out(87),
            data_re_out(6) => data_re_out(103),
            data_re_out(7) => data_re_out(119),
            data_re_out(8) => data_re_out(135),
            data_re_out(9) => data_re_out(151),
            data_re_out(10) => data_re_out(167),
            data_re_out(11) => data_re_out(183),
            data_re_out(12) => data_re_out(199),
            data_re_out(13) => data_re_out(215),
            data_re_out(14) => data_re_out(231),
            data_re_out(15) => data_re_out(247),
            data_re_out(16) => data_re_out(263),
            data_re_out(17) => data_re_out(279),
            data_re_out(18) => data_re_out(295),
            data_re_out(19) => data_re_out(311),
            data_re_out(20) => data_re_out(327),
            data_re_out(21) => data_re_out(343),
            data_re_out(22) => data_re_out(359),
            data_re_out(23) => data_re_out(375),
            data_re_out(24) => data_re_out(391),
            data_re_out(25) => data_re_out(407),
            data_re_out(26) => data_re_out(423),
            data_re_out(27) => data_re_out(439),
            data_re_out(28) => data_re_out(455),
            data_re_out(29) => data_re_out(471),
            data_re_out(30) => data_re_out(487),
            data_re_out(31) => data_re_out(503),
            data_im_out(0) => data_im_out(7),
            data_im_out(1) => data_im_out(23),
            data_im_out(2) => data_im_out(39),
            data_im_out(3) => data_im_out(55),
            data_im_out(4) => data_im_out(71),
            data_im_out(5) => data_im_out(87),
            data_im_out(6) => data_im_out(103),
            data_im_out(7) => data_im_out(119),
            data_im_out(8) => data_im_out(135),
            data_im_out(9) => data_im_out(151),
            data_im_out(10) => data_im_out(167),
            data_im_out(11) => data_im_out(183),
            data_im_out(12) => data_im_out(199),
            data_im_out(13) => data_im_out(215),
            data_im_out(14) => data_im_out(231),
            data_im_out(15) => data_im_out(247),
            data_im_out(16) => data_im_out(263),
            data_im_out(17) => data_im_out(279),
            data_im_out(18) => data_im_out(295),
            data_im_out(19) => data_im_out(311),
            data_im_out(20) => data_im_out(327),
            data_im_out(21) => data_im_out(343),
            data_im_out(22) => data_im_out(359),
            data_im_out(23) => data_im_out(375),
            data_im_out(24) => data_im_out(391),
            data_im_out(25) => data_im_out(407),
            data_im_out(26) => data_im_out(423),
            data_im_out(27) => data_im_out(439),
            data_im_out(28) => data_im_out(455),
            data_im_out(29) => data_im_out(471),
            data_im_out(30) => data_im_out(487),
            data_im_out(31) => data_im_out(503)
        );           

    URFFT_PT32_8 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(256),
            data_re_in(1) => mul_re_out(257),
            data_re_in(2) => mul_re_out(258),
            data_re_in(3) => mul_re_out(259),
            data_re_in(4) => mul_re_out(260),
            data_re_in(5) => mul_re_out(261),
            data_re_in(6) => mul_re_out(262),
            data_re_in(7) => mul_re_out(263),
            data_re_in(8) => mul_re_out(264),
            data_re_in(9) => mul_re_out(265),
            data_re_in(10) => mul_re_out(266),
            data_re_in(11) => mul_re_out(267),
            data_re_in(12) => mul_re_out(268),
            data_re_in(13) => mul_re_out(269),
            data_re_in(14) => mul_re_out(270),
            data_re_in(15) => mul_re_out(271),
            data_re_in(16) => mul_re_out(272),
            data_re_in(17) => mul_re_out(273),
            data_re_in(18) => mul_re_out(274),
            data_re_in(19) => mul_re_out(275),
            data_re_in(20) => mul_re_out(276),
            data_re_in(21) => mul_re_out(277),
            data_re_in(22) => mul_re_out(278),
            data_re_in(23) => mul_re_out(279),
            data_re_in(24) => mul_re_out(280),
            data_re_in(25) => mul_re_out(281),
            data_re_in(26) => mul_re_out(282),
            data_re_in(27) => mul_re_out(283),
            data_re_in(28) => mul_re_out(284),
            data_re_in(29) => mul_re_out(285),
            data_re_in(30) => mul_re_out(286),
            data_re_in(31) => mul_re_out(287),
            data_im_in(0) => mul_im_out(256),
            data_im_in(1) => mul_im_out(257),
            data_im_in(2) => mul_im_out(258),
            data_im_in(3) => mul_im_out(259),
            data_im_in(4) => mul_im_out(260),
            data_im_in(5) => mul_im_out(261),
            data_im_in(6) => mul_im_out(262),
            data_im_in(7) => mul_im_out(263),
            data_im_in(8) => mul_im_out(264),
            data_im_in(9) => mul_im_out(265),
            data_im_in(10) => mul_im_out(266),
            data_im_in(11) => mul_im_out(267),
            data_im_in(12) => mul_im_out(268),
            data_im_in(13) => mul_im_out(269),
            data_im_in(14) => mul_im_out(270),
            data_im_in(15) => mul_im_out(271),
            data_im_in(16) => mul_im_out(272),
            data_im_in(17) => mul_im_out(273),
            data_im_in(18) => mul_im_out(274),
            data_im_in(19) => mul_im_out(275),
            data_im_in(20) => mul_im_out(276),
            data_im_in(21) => mul_im_out(277),
            data_im_in(22) => mul_im_out(278),
            data_im_in(23) => mul_im_out(279),
            data_im_in(24) => mul_im_out(280),
            data_im_in(25) => mul_im_out(281),
            data_im_in(26) => mul_im_out(282),
            data_im_in(27) => mul_im_out(283),
            data_im_in(28) => mul_im_out(284),
            data_im_in(29) => mul_im_out(285),
            data_im_in(30) => mul_im_out(286),
            data_im_in(31) => mul_im_out(287),
            data_re_out(0) => data_re_out(8),
            data_re_out(1) => data_re_out(24),
            data_re_out(2) => data_re_out(40),
            data_re_out(3) => data_re_out(56),
            data_re_out(4) => data_re_out(72),
            data_re_out(5) => data_re_out(88),
            data_re_out(6) => data_re_out(104),
            data_re_out(7) => data_re_out(120),
            data_re_out(8) => data_re_out(136),
            data_re_out(9) => data_re_out(152),
            data_re_out(10) => data_re_out(168),
            data_re_out(11) => data_re_out(184),
            data_re_out(12) => data_re_out(200),
            data_re_out(13) => data_re_out(216),
            data_re_out(14) => data_re_out(232),
            data_re_out(15) => data_re_out(248),
            data_re_out(16) => data_re_out(264),
            data_re_out(17) => data_re_out(280),
            data_re_out(18) => data_re_out(296),
            data_re_out(19) => data_re_out(312),
            data_re_out(20) => data_re_out(328),
            data_re_out(21) => data_re_out(344),
            data_re_out(22) => data_re_out(360),
            data_re_out(23) => data_re_out(376),
            data_re_out(24) => data_re_out(392),
            data_re_out(25) => data_re_out(408),
            data_re_out(26) => data_re_out(424),
            data_re_out(27) => data_re_out(440),
            data_re_out(28) => data_re_out(456),
            data_re_out(29) => data_re_out(472),
            data_re_out(30) => data_re_out(488),
            data_re_out(31) => data_re_out(504),
            data_im_out(0) => data_im_out(8),
            data_im_out(1) => data_im_out(24),
            data_im_out(2) => data_im_out(40),
            data_im_out(3) => data_im_out(56),
            data_im_out(4) => data_im_out(72),
            data_im_out(5) => data_im_out(88),
            data_im_out(6) => data_im_out(104),
            data_im_out(7) => data_im_out(120),
            data_im_out(8) => data_im_out(136),
            data_im_out(9) => data_im_out(152),
            data_im_out(10) => data_im_out(168),
            data_im_out(11) => data_im_out(184),
            data_im_out(12) => data_im_out(200),
            data_im_out(13) => data_im_out(216),
            data_im_out(14) => data_im_out(232),
            data_im_out(15) => data_im_out(248),
            data_im_out(16) => data_im_out(264),
            data_im_out(17) => data_im_out(280),
            data_im_out(18) => data_im_out(296),
            data_im_out(19) => data_im_out(312),
            data_im_out(20) => data_im_out(328),
            data_im_out(21) => data_im_out(344),
            data_im_out(22) => data_im_out(360),
            data_im_out(23) => data_im_out(376),
            data_im_out(24) => data_im_out(392),
            data_im_out(25) => data_im_out(408),
            data_im_out(26) => data_im_out(424),
            data_im_out(27) => data_im_out(440),
            data_im_out(28) => data_im_out(456),
            data_im_out(29) => data_im_out(472),
            data_im_out(30) => data_im_out(488),
            data_im_out(31) => data_im_out(504)
        );           

    URFFT_PT32_9 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(288),
            data_re_in(1) => mul_re_out(289),
            data_re_in(2) => mul_re_out(290),
            data_re_in(3) => mul_re_out(291),
            data_re_in(4) => mul_re_out(292),
            data_re_in(5) => mul_re_out(293),
            data_re_in(6) => mul_re_out(294),
            data_re_in(7) => mul_re_out(295),
            data_re_in(8) => mul_re_out(296),
            data_re_in(9) => mul_re_out(297),
            data_re_in(10) => mul_re_out(298),
            data_re_in(11) => mul_re_out(299),
            data_re_in(12) => mul_re_out(300),
            data_re_in(13) => mul_re_out(301),
            data_re_in(14) => mul_re_out(302),
            data_re_in(15) => mul_re_out(303),
            data_re_in(16) => mul_re_out(304),
            data_re_in(17) => mul_re_out(305),
            data_re_in(18) => mul_re_out(306),
            data_re_in(19) => mul_re_out(307),
            data_re_in(20) => mul_re_out(308),
            data_re_in(21) => mul_re_out(309),
            data_re_in(22) => mul_re_out(310),
            data_re_in(23) => mul_re_out(311),
            data_re_in(24) => mul_re_out(312),
            data_re_in(25) => mul_re_out(313),
            data_re_in(26) => mul_re_out(314),
            data_re_in(27) => mul_re_out(315),
            data_re_in(28) => mul_re_out(316),
            data_re_in(29) => mul_re_out(317),
            data_re_in(30) => mul_re_out(318),
            data_re_in(31) => mul_re_out(319),
            data_im_in(0) => mul_im_out(288),
            data_im_in(1) => mul_im_out(289),
            data_im_in(2) => mul_im_out(290),
            data_im_in(3) => mul_im_out(291),
            data_im_in(4) => mul_im_out(292),
            data_im_in(5) => mul_im_out(293),
            data_im_in(6) => mul_im_out(294),
            data_im_in(7) => mul_im_out(295),
            data_im_in(8) => mul_im_out(296),
            data_im_in(9) => mul_im_out(297),
            data_im_in(10) => mul_im_out(298),
            data_im_in(11) => mul_im_out(299),
            data_im_in(12) => mul_im_out(300),
            data_im_in(13) => mul_im_out(301),
            data_im_in(14) => mul_im_out(302),
            data_im_in(15) => mul_im_out(303),
            data_im_in(16) => mul_im_out(304),
            data_im_in(17) => mul_im_out(305),
            data_im_in(18) => mul_im_out(306),
            data_im_in(19) => mul_im_out(307),
            data_im_in(20) => mul_im_out(308),
            data_im_in(21) => mul_im_out(309),
            data_im_in(22) => mul_im_out(310),
            data_im_in(23) => mul_im_out(311),
            data_im_in(24) => mul_im_out(312),
            data_im_in(25) => mul_im_out(313),
            data_im_in(26) => mul_im_out(314),
            data_im_in(27) => mul_im_out(315),
            data_im_in(28) => mul_im_out(316),
            data_im_in(29) => mul_im_out(317),
            data_im_in(30) => mul_im_out(318),
            data_im_in(31) => mul_im_out(319),
            data_re_out(0) => data_re_out(9),
            data_re_out(1) => data_re_out(25),
            data_re_out(2) => data_re_out(41),
            data_re_out(3) => data_re_out(57),
            data_re_out(4) => data_re_out(73),
            data_re_out(5) => data_re_out(89),
            data_re_out(6) => data_re_out(105),
            data_re_out(7) => data_re_out(121),
            data_re_out(8) => data_re_out(137),
            data_re_out(9) => data_re_out(153),
            data_re_out(10) => data_re_out(169),
            data_re_out(11) => data_re_out(185),
            data_re_out(12) => data_re_out(201),
            data_re_out(13) => data_re_out(217),
            data_re_out(14) => data_re_out(233),
            data_re_out(15) => data_re_out(249),
            data_re_out(16) => data_re_out(265),
            data_re_out(17) => data_re_out(281),
            data_re_out(18) => data_re_out(297),
            data_re_out(19) => data_re_out(313),
            data_re_out(20) => data_re_out(329),
            data_re_out(21) => data_re_out(345),
            data_re_out(22) => data_re_out(361),
            data_re_out(23) => data_re_out(377),
            data_re_out(24) => data_re_out(393),
            data_re_out(25) => data_re_out(409),
            data_re_out(26) => data_re_out(425),
            data_re_out(27) => data_re_out(441),
            data_re_out(28) => data_re_out(457),
            data_re_out(29) => data_re_out(473),
            data_re_out(30) => data_re_out(489),
            data_re_out(31) => data_re_out(505),
            data_im_out(0) => data_im_out(9),
            data_im_out(1) => data_im_out(25),
            data_im_out(2) => data_im_out(41),
            data_im_out(3) => data_im_out(57),
            data_im_out(4) => data_im_out(73),
            data_im_out(5) => data_im_out(89),
            data_im_out(6) => data_im_out(105),
            data_im_out(7) => data_im_out(121),
            data_im_out(8) => data_im_out(137),
            data_im_out(9) => data_im_out(153),
            data_im_out(10) => data_im_out(169),
            data_im_out(11) => data_im_out(185),
            data_im_out(12) => data_im_out(201),
            data_im_out(13) => data_im_out(217),
            data_im_out(14) => data_im_out(233),
            data_im_out(15) => data_im_out(249),
            data_im_out(16) => data_im_out(265),
            data_im_out(17) => data_im_out(281),
            data_im_out(18) => data_im_out(297),
            data_im_out(19) => data_im_out(313),
            data_im_out(20) => data_im_out(329),
            data_im_out(21) => data_im_out(345),
            data_im_out(22) => data_im_out(361),
            data_im_out(23) => data_im_out(377),
            data_im_out(24) => data_im_out(393),
            data_im_out(25) => data_im_out(409),
            data_im_out(26) => data_im_out(425),
            data_im_out(27) => data_im_out(441),
            data_im_out(28) => data_im_out(457),
            data_im_out(29) => data_im_out(473),
            data_im_out(30) => data_im_out(489),
            data_im_out(31) => data_im_out(505)
        );           

    URFFT_PT32_10 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(320),
            data_re_in(1) => mul_re_out(321),
            data_re_in(2) => mul_re_out(322),
            data_re_in(3) => mul_re_out(323),
            data_re_in(4) => mul_re_out(324),
            data_re_in(5) => mul_re_out(325),
            data_re_in(6) => mul_re_out(326),
            data_re_in(7) => mul_re_out(327),
            data_re_in(8) => mul_re_out(328),
            data_re_in(9) => mul_re_out(329),
            data_re_in(10) => mul_re_out(330),
            data_re_in(11) => mul_re_out(331),
            data_re_in(12) => mul_re_out(332),
            data_re_in(13) => mul_re_out(333),
            data_re_in(14) => mul_re_out(334),
            data_re_in(15) => mul_re_out(335),
            data_re_in(16) => mul_re_out(336),
            data_re_in(17) => mul_re_out(337),
            data_re_in(18) => mul_re_out(338),
            data_re_in(19) => mul_re_out(339),
            data_re_in(20) => mul_re_out(340),
            data_re_in(21) => mul_re_out(341),
            data_re_in(22) => mul_re_out(342),
            data_re_in(23) => mul_re_out(343),
            data_re_in(24) => mul_re_out(344),
            data_re_in(25) => mul_re_out(345),
            data_re_in(26) => mul_re_out(346),
            data_re_in(27) => mul_re_out(347),
            data_re_in(28) => mul_re_out(348),
            data_re_in(29) => mul_re_out(349),
            data_re_in(30) => mul_re_out(350),
            data_re_in(31) => mul_re_out(351),
            data_im_in(0) => mul_im_out(320),
            data_im_in(1) => mul_im_out(321),
            data_im_in(2) => mul_im_out(322),
            data_im_in(3) => mul_im_out(323),
            data_im_in(4) => mul_im_out(324),
            data_im_in(5) => mul_im_out(325),
            data_im_in(6) => mul_im_out(326),
            data_im_in(7) => mul_im_out(327),
            data_im_in(8) => mul_im_out(328),
            data_im_in(9) => mul_im_out(329),
            data_im_in(10) => mul_im_out(330),
            data_im_in(11) => mul_im_out(331),
            data_im_in(12) => mul_im_out(332),
            data_im_in(13) => mul_im_out(333),
            data_im_in(14) => mul_im_out(334),
            data_im_in(15) => mul_im_out(335),
            data_im_in(16) => mul_im_out(336),
            data_im_in(17) => mul_im_out(337),
            data_im_in(18) => mul_im_out(338),
            data_im_in(19) => mul_im_out(339),
            data_im_in(20) => mul_im_out(340),
            data_im_in(21) => mul_im_out(341),
            data_im_in(22) => mul_im_out(342),
            data_im_in(23) => mul_im_out(343),
            data_im_in(24) => mul_im_out(344),
            data_im_in(25) => mul_im_out(345),
            data_im_in(26) => mul_im_out(346),
            data_im_in(27) => mul_im_out(347),
            data_im_in(28) => mul_im_out(348),
            data_im_in(29) => mul_im_out(349),
            data_im_in(30) => mul_im_out(350),
            data_im_in(31) => mul_im_out(351),
            data_re_out(0) => data_re_out(10),
            data_re_out(1) => data_re_out(26),
            data_re_out(2) => data_re_out(42),
            data_re_out(3) => data_re_out(58),
            data_re_out(4) => data_re_out(74),
            data_re_out(5) => data_re_out(90),
            data_re_out(6) => data_re_out(106),
            data_re_out(7) => data_re_out(122),
            data_re_out(8) => data_re_out(138),
            data_re_out(9) => data_re_out(154),
            data_re_out(10) => data_re_out(170),
            data_re_out(11) => data_re_out(186),
            data_re_out(12) => data_re_out(202),
            data_re_out(13) => data_re_out(218),
            data_re_out(14) => data_re_out(234),
            data_re_out(15) => data_re_out(250),
            data_re_out(16) => data_re_out(266),
            data_re_out(17) => data_re_out(282),
            data_re_out(18) => data_re_out(298),
            data_re_out(19) => data_re_out(314),
            data_re_out(20) => data_re_out(330),
            data_re_out(21) => data_re_out(346),
            data_re_out(22) => data_re_out(362),
            data_re_out(23) => data_re_out(378),
            data_re_out(24) => data_re_out(394),
            data_re_out(25) => data_re_out(410),
            data_re_out(26) => data_re_out(426),
            data_re_out(27) => data_re_out(442),
            data_re_out(28) => data_re_out(458),
            data_re_out(29) => data_re_out(474),
            data_re_out(30) => data_re_out(490),
            data_re_out(31) => data_re_out(506),
            data_im_out(0) => data_im_out(10),
            data_im_out(1) => data_im_out(26),
            data_im_out(2) => data_im_out(42),
            data_im_out(3) => data_im_out(58),
            data_im_out(4) => data_im_out(74),
            data_im_out(5) => data_im_out(90),
            data_im_out(6) => data_im_out(106),
            data_im_out(7) => data_im_out(122),
            data_im_out(8) => data_im_out(138),
            data_im_out(9) => data_im_out(154),
            data_im_out(10) => data_im_out(170),
            data_im_out(11) => data_im_out(186),
            data_im_out(12) => data_im_out(202),
            data_im_out(13) => data_im_out(218),
            data_im_out(14) => data_im_out(234),
            data_im_out(15) => data_im_out(250),
            data_im_out(16) => data_im_out(266),
            data_im_out(17) => data_im_out(282),
            data_im_out(18) => data_im_out(298),
            data_im_out(19) => data_im_out(314),
            data_im_out(20) => data_im_out(330),
            data_im_out(21) => data_im_out(346),
            data_im_out(22) => data_im_out(362),
            data_im_out(23) => data_im_out(378),
            data_im_out(24) => data_im_out(394),
            data_im_out(25) => data_im_out(410),
            data_im_out(26) => data_im_out(426),
            data_im_out(27) => data_im_out(442),
            data_im_out(28) => data_im_out(458),
            data_im_out(29) => data_im_out(474),
            data_im_out(30) => data_im_out(490),
            data_im_out(31) => data_im_out(506)
        );           

    URFFT_PT32_11 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(352),
            data_re_in(1) => mul_re_out(353),
            data_re_in(2) => mul_re_out(354),
            data_re_in(3) => mul_re_out(355),
            data_re_in(4) => mul_re_out(356),
            data_re_in(5) => mul_re_out(357),
            data_re_in(6) => mul_re_out(358),
            data_re_in(7) => mul_re_out(359),
            data_re_in(8) => mul_re_out(360),
            data_re_in(9) => mul_re_out(361),
            data_re_in(10) => mul_re_out(362),
            data_re_in(11) => mul_re_out(363),
            data_re_in(12) => mul_re_out(364),
            data_re_in(13) => mul_re_out(365),
            data_re_in(14) => mul_re_out(366),
            data_re_in(15) => mul_re_out(367),
            data_re_in(16) => mul_re_out(368),
            data_re_in(17) => mul_re_out(369),
            data_re_in(18) => mul_re_out(370),
            data_re_in(19) => mul_re_out(371),
            data_re_in(20) => mul_re_out(372),
            data_re_in(21) => mul_re_out(373),
            data_re_in(22) => mul_re_out(374),
            data_re_in(23) => mul_re_out(375),
            data_re_in(24) => mul_re_out(376),
            data_re_in(25) => mul_re_out(377),
            data_re_in(26) => mul_re_out(378),
            data_re_in(27) => mul_re_out(379),
            data_re_in(28) => mul_re_out(380),
            data_re_in(29) => mul_re_out(381),
            data_re_in(30) => mul_re_out(382),
            data_re_in(31) => mul_re_out(383),
            data_im_in(0) => mul_im_out(352),
            data_im_in(1) => mul_im_out(353),
            data_im_in(2) => mul_im_out(354),
            data_im_in(3) => mul_im_out(355),
            data_im_in(4) => mul_im_out(356),
            data_im_in(5) => mul_im_out(357),
            data_im_in(6) => mul_im_out(358),
            data_im_in(7) => mul_im_out(359),
            data_im_in(8) => mul_im_out(360),
            data_im_in(9) => mul_im_out(361),
            data_im_in(10) => mul_im_out(362),
            data_im_in(11) => mul_im_out(363),
            data_im_in(12) => mul_im_out(364),
            data_im_in(13) => mul_im_out(365),
            data_im_in(14) => mul_im_out(366),
            data_im_in(15) => mul_im_out(367),
            data_im_in(16) => mul_im_out(368),
            data_im_in(17) => mul_im_out(369),
            data_im_in(18) => mul_im_out(370),
            data_im_in(19) => mul_im_out(371),
            data_im_in(20) => mul_im_out(372),
            data_im_in(21) => mul_im_out(373),
            data_im_in(22) => mul_im_out(374),
            data_im_in(23) => mul_im_out(375),
            data_im_in(24) => mul_im_out(376),
            data_im_in(25) => mul_im_out(377),
            data_im_in(26) => mul_im_out(378),
            data_im_in(27) => mul_im_out(379),
            data_im_in(28) => mul_im_out(380),
            data_im_in(29) => mul_im_out(381),
            data_im_in(30) => mul_im_out(382),
            data_im_in(31) => mul_im_out(383),
            data_re_out(0) => data_re_out(11),
            data_re_out(1) => data_re_out(27),
            data_re_out(2) => data_re_out(43),
            data_re_out(3) => data_re_out(59),
            data_re_out(4) => data_re_out(75),
            data_re_out(5) => data_re_out(91),
            data_re_out(6) => data_re_out(107),
            data_re_out(7) => data_re_out(123),
            data_re_out(8) => data_re_out(139),
            data_re_out(9) => data_re_out(155),
            data_re_out(10) => data_re_out(171),
            data_re_out(11) => data_re_out(187),
            data_re_out(12) => data_re_out(203),
            data_re_out(13) => data_re_out(219),
            data_re_out(14) => data_re_out(235),
            data_re_out(15) => data_re_out(251),
            data_re_out(16) => data_re_out(267),
            data_re_out(17) => data_re_out(283),
            data_re_out(18) => data_re_out(299),
            data_re_out(19) => data_re_out(315),
            data_re_out(20) => data_re_out(331),
            data_re_out(21) => data_re_out(347),
            data_re_out(22) => data_re_out(363),
            data_re_out(23) => data_re_out(379),
            data_re_out(24) => data_re_out(395),
            data_re_out(25) => data_re_out(411),
            data_re_out(26) => data_re_out(427),
            data_re_out(27) => data_re_out(443),
            data_re_out(28) => data_re_out(459),
            data_re_out(29) => data_re_out(475),
            data_re_out(30) => data_re_out(491),
            data_re_out(31) => data_re_out(507),
            data_im_out(0) => data_im_out(11),
            data_im_out(1) => data_im_out(27),
            data_im_out(2) => data_im_out(43),
            data_im_out(3) => data_im_out(59),
            data_im_out(4) => data_im_out(75),
            data_im_out(5) => data_im_out(91),
            data_im_out(6) => data_im_out(107),
            data_im_out(7) => data_im_out(123),
            data_im_out(8) => data_im_out(139),
            data_im_out(9) => data_im_out(155),
            data_im_out(10) => data_im_out(171),
            data_im_out(11) => data_im_out(187),
            data_im_out(12) => data_im_out(203),
            data_im_out(13) => data_im_out(219),
            data_im_out(14) => data_im_out(235),
            data_im_out(15) => data_im_out(251),
            data_im_out(16) => data_im_out(267),
            data_im_out(17) => data_im_out(283),
            data_im_out(18) => data_im_out(299),
            data_im_out(19) => data_im_out(315),
            data_im_out(20) => data_im_out(331),
            data_im_out(21) => data_im_out(347),
            data_im_out(22) => data_im_out(363),
            data_im_out(23) => data_im_out(379),
            data_im_out(24) => data_im_out(395),
            data_im_out(25) => data_im_out(411),
            data_im_out(26) => data_im_out(427),
            data_im_out(27) => data_im_out(443),
            data_im_out(28) => data_im_out(459),
            data_im_out(29) => data_im_out(475),
            data_im_out(30) => data_im_out(491),
            data_im_out(31) => data_im_out(507)
        );           

    URFFT_PT32_12 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(384),
            data_re_in(1) => mul_re_out(385),
            data_re_in(2) => mul_re_out(386),
            data_re_in(3) => mul_re_out(387),
            data_re_in(4) => mul_re_out(388),
            data_re_in(5) => mul_re_out(389),
            data_re_in(6) => mul_re_out(390),
            data_re_in(7) => mul_re_out(391),
            data_re_in(8) => mul_re_out(392),
            data_re_in(9) => mul_re_out(393),
            data_re_in(10) => mul_re_out(394),
            data_re_in(11) => mul_re_out(395),
            data_re_in(12) => mul_re_out(396),
            data_re_in(13) => mul_re_out(397),
            data_re_in(14) => mul_re_out(398),
            data_re_in(15) => mul_re_out(399),
            data_re_in(16) => mul_re_out(400),
            data_re_in(17) => mul_re_out(401),
            data_re_in(18) => mul_re_out(402),
            data_re_in(19) => mul_re_out(403),
            data_re_in(20) => mul_re_out(404),
            data_re_in(21) => mul_re_out(405),
            data_re_in(22) => mul_re_out(406),
            data_re_in(23) => mul_re_out(407),
            data_re_in(24) => mul_re_out(408),
            data_re_in(25) => mul_re_out(409),
            data_re_in(26) => mul_re_out(410),
            data_re_in(27) => mul_re_out(411),
            data_re_in(28) => mul_re_out(412),
            data_re_in(29) => mul_re_out(413),
            data_re_in(30) => mul_re_out(414),
            data_re_in(31) => mul_re_out(415),
            data_im_in(0) => mul_im_out(384),
            data_im_in(1) => mul_im_out(385),
            data_im_in(2) => mul_im_out(386),
            data_im_in(3) => mul_im_out(387),
            data_im_in(4) => mul_im_out(388),
            data_im_in(5) => mul_im_out(389),
            data_im_in(6) => mul_im_out(390),
            data_im_in(7) => mul_im_out(391),
            data_im_in(8) => mul_im_out(392),
            data_im_in(9) => mul_im_out(393),
            data_im_in(10) => mul_im_out(394),
            data_im_in(11) => mul_im_out(395),
            data_im_in(12) => mul_im_out(396),
            data_im_in(13) => mul_im_out(397),
            data_im_in(14) => mul_im_out(398),
            data_im_in(15) => mul_im_out(399),
            data_im_in(16) => mul_im_out(400),
            data_im_in(17) => mul_im_out(401),
            data_im_in(18) => mul_im_out(402),
            data_im_in(19) => mul_im_out(403),
            data_im_in(20) => mul_im_out(404),
            data_im_in(21) => mul_im_out(405),
            data_im_in(22) => mul_im_out(406),
            data_im_in(23) => mul_im_out(407),
            data_im_in(24) => mul_im_out(408),
            data_im_in(25) => mul_im_out(409),
            data_im_in(26) => mul_im_out(410),
            data_im_in(27) => mul_im_out(411),
            data_im_in(28) => mul_im_out(412),
            data_im_in(29) => mul_im_out(413),
            data_im_in(30) => mul_im_out(414),
            data_im_in(31) => mul_im_out(415),
            data_re_out(0) => data_re_out(12),
            data_re_out(1) => data_re_out(28),
            data_re_out(2) => data_re_out(44),
            data_re_out(3) => data_re_out(60),
            data_re_out(4) => data_re_out(76),
            data_re_out(5) => data_re_out(92),
            data_re_out(6) => data_re_out(108),
            data_re_out(7) => data_re_out(124),
            data_re_out(8) => data_re_out(140),
            data_re_out(9) => data_re_out(156),
            data_re_out(10) => data_re_out(172),
            data_re_out(11) => data_re_out(188),
            data_re_out(12) => data_re_out(204),
            data_re_out(13) => data_re_out(220),
            data_re_out(14) => data_re_out(236),
            data_re_out(15) => data_re_out(252),
            data_re_out(16) => data_re_out(268),
            data_re_out(17) => data_re_out(284),
            data_re_out(18) => data_re_out(300),
            data_re_out(19) => data_re_out(316),
            data_re_out(20) => data_re_out(332),
            data_re_out(21) => data_re_out(348),
            data_re_out(22) => data_re_out(364),
            data_re_out(23) => data_re_out(380),
            data_re_out(24) => data_re_out(396),
            data_re_out(25) => data_re_out(412),
            data_re_out(26) => data_re_out(428),
            data_re_out(27) => data_re_out(444),
            data_re_out(28) => data_re_out(460),
            data_re_out(29) => data_re_out(476),
            data_re_out(30) => data_re_out(492),
            data_re_out(31) => data_re_out(508),
            data_im_out(0) => data_im_out(12),
            data_im_out(1) => data_im_out(28),
            data_im_out(2) => data_im_out(44),
            data_im_out(3) => data_im_out(60),
            data_im_out(4) => data_im_out(76),
            data_im_out(5) => data_im_out(92),
            data_im_out(6) => data_im_out(108),
            data_im_out(7) => data_im_out(124),
            data_im_out(8) => data_im_out(140),
            data_im_out(9) => data_im_out(156),
            data_im_out(10) => data_im_out(172),
            data_im_out(11) => data_im_out(188),
            data_im_out(12) => data_im_out(204),
            data_im_out(13) => data_im_out(220),
            data_im_out(14) => data_im_out(236),
            data_im_out(15) => data_im_out(252),
            data_im_out(16) => data_im_out(268),
            data_im_out(17) => data_im_out(284),
            data_im_out(18) => data_im_out(300),
            data_im_out(19) => data_im_out(316),
            data_im_out(20) => data_im_out(332),
            data_im_out(21) => data_im_out(348),
            data_im_out(22) => data_im_out(364),
            data_im_out(23) => data_im_out(380),
            data_im_out(24) => data_im_out(396),
            data_im_out(25) => data_im_out(412),
            data_im_out(26) => data_im_out(428),
            data_im_out(27) => data_im_out(444),
            data_im_out(28) => data_im_out(460),
            data_im_out(29) => data_im_out(476),
            data_im_out(30) => data_im_out(492),
            data_im_out(31) => data_im_out(508)
        );           

    URFFT_PT32_13 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(416),
            data_re_in(1) => mul_re_out(417),
            data_re_in(2) => mul_re_out(418),
            data_re_in(3) => mul_re_out(419),
            data_re_in(4) => mul_re_out(420),
            data_re_in(5) => mul_re_out(421),
            data_re_in(6) => mul_re_out(422),
            data_re_in(7) => mul_re_out(423),
            data_re_in(8) => mul_re_out(424),
            data_re_in(9) => mul_re_out(425),
            data_re_in(10) => mul_re_out(426),
            data_re_in(11) => mul_re_out(427),
            data_re_in(12) => mul_re_out(428),
            data_re_in(13) => mul_re_out(429),
            data_re_in(14) => mul_re_out(430),
            data_re_in(15) => mul_re_out(431),
            data_re_in(16) => mul_re_out(432),
            data_re_in(17) => mul_re_out(433),
            data_re_in(18) => mul_re_out(434),
            data_re_in(19) => mul_re_out(435),
            data_re_in(20) => mul_re_out(436),
            data_re_in(21) => mul_re_out(437),
            data_re_in(22) => mul_re_out(438),
            data_re_in(23) => mul_re_out(439),
            data_re_in(24) => mul_re_out(440),
            data_re_in(25) => mul_re_out(441),
            data_re_in(26) => mul_re_out(442),
            data_re_in(27) => mul_re_out(443),
            data_re_in(28) => mul_re_out(444),
            data_re_in(29) => mul_re_out(445),
            data_re_in(30) => mul_re_out(446),
            data_re_in(31) => mul_re_out(447),
            data_im_in(0) => mul_im_out(416),
            data_im_in(1) => mul_im_out(417),
            data_im_in(2) => mul_im_out(418),
            data_im_in(3) => mul_im_out(419),
            data_im_in(4) => mul_im_out(420),
            data_im_in(5) => mul_im_out(421),
            data_im_in(6) => mul_im_out(422),
            data_im_in(7) => mul_im_out(423),
            data_im_in(8) => mul_im_out(424),
            data_im_in(9) => mul_im_out(425),
            data_im_in(10) => mul_im_out(426),
            data_im_in(11) => mul_im_out(427),
            data_im_in(12) => mul_im_out(428),
            data_im_in(13) => mul_im_out(429),
            data_im_in(14) => mul_im_out(430),
            data_im_in(15) => mul_im_out(431),
            data_im_in(16) => mul_im_out(432),
            data_im_in(17) => mul_im_out(433),
            data_im_in(18) => mul_im_out(434),
            data_im_in(19) => mul_im_out(435),
            data_im_in(20) => mul_im_out(436),
            data_im_in(21) => mul_im_out(437),
            data_im_in(22) => mul_im_out(438),
            data_im_in(23) => mul_im_out(439),
            data_im_in(24) => mul_im_out(440),
            data_im_in(25) => mul_im_out(441),
            data_im_in(26) => mul_im_out(442),
            data_im_in(27) => mul_im_out(443),
            data_im_in(28) => mul_im_out(444),
            data_im_in(29) => mul_im_out(445),
            data_im_in(30) => mul_im_out(446),
            data_im_in(31) => mul_im_out(447),
            data_re_out(0) => data_re_out(13),
            data_re_out(1) => data_re_out(29),
            data_re_out(2) => data_re_out(45),
            data_re_out(3) => data_re_out(61),
            data_re_out(4) => data_re_out(77),
            data_re_out(5) => data_re_out(93),
            data_re_out(6) => data_re_out(109),
            data_re_out(7) => data_re_out(125),
            data_re_out(8) => data_re_out(141),
            data_re_out(9) => data_re_out(157),
            data_re_out(10) => data_re_out(173),
            data_re_out(11) => data_re_out(189),
            data_re_out(12) => data_re_out(205),
            data_re_out(13) => data_re_out(221),
            data_re_out(14) => data_re_out(237),
            data_re_out(15) => data_re_out(253),
            data_re_out(16) => data_re_out(269),
            data_re_out(17) => data_re_out(285),
            data_re_out(18) => data_re_out(301),
            data_re_out(19) => data_re_out(317),
            data_re_out(20) => data_re_out(333),
            data_re_out(21) => data_re_out(349),
            data_re_out(22) => data_re_out(365),
            data_re_out(23) => data_re_out(381),
            data_re_out(24) => data_re_out(397),
            data_re_out(25) => data_re_out(413),
            data_re_out(26) => data_re_out(429),
            data_re_out(27) => data_re_out(445),
            data_re_out(28) => data_re_out(461),
            data_re_out(29) => data_re_out(477),
            data_re_out(30) => data_re_out(493),
            data_re_out(31) => data_re_out(509),
            data_im_out(0) => data_im_out(13),
            data_im_out(1) => data_im_out(29),
            data_im_out(2) => data_im_out(45),
            data_im_out(3) => data_im_out(61),
            data_im_out(4) => data_im_out(77),
            data_im_out(5) => data_im_out(93),
            data_im_out(6) => data_im_out(109),
            data_im_out(7) => data_im_out(125),
            data_im_out(8) => data_im_out(141),
            data_im_out(9) => data_im_out(157),
            data_im_out(10) => data_im_out(173),
            data_im_out(11) => data_im_out(189),
            data_im_out(12) => data_im_out(205),
            data_im_out(13) => data_im_out(221),
            data_im_out(14) => data_im_out(237),
            data_im_out(15) => data_im_out(253),
            data_im_out(16) => data_im_out(269),
            data_im_out(17) => data_im_out(285),
            data_im_out(18) => data_im_out(301),
            data_im_out(19) => data_im_out(317),
            data_im_out(20) => data_im_out(333),
            data_im_out(21) => data_im_out(349),
            data_im_out(22) => data_im_out(365),
            data_im_out(23) => data_im_out(381),
            data_im_out(24) => data_im_out(397),
            data_im_out(25) => data_im_out(413),
            data_im_out(26) => data_im_out(429),
            data_im_out(27) => data_im_out(445),
            data_im_out(28) => data_im_out(461),
            data_im_out(29) => data_im_out(477),
            data_im_out(30) => data_im_out(493),
            data_im_out(31) => data_im_out(509)
        );           

    URFFT_PT32_14 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(448),
            data_re_in(1) => mul_re_out(449),
            data_re_in(2) => mul_re_out(450),
            data_re_in(3) => mul_re_out(451),
            data_re_in(4) => mul_re_out(452),
            data_re_in(5) => mul_re_out(453),
            data_re_in(6) => mul_re_out(454),
            data_re_in(7) => mul_re_out(455),
            data_re_in(8) => mul_re_out(456),
            data_re_in(9) => mul_re_out(457),
            data_re_in(10) => mul_re_out(458),
            data_re_in(11) => mul_re_out(459),
            data_re_in(12) => mul_re_out(460),
            data_re_in(13) => mul_re_out(461),
            data_re_in(14) => mul_re_out(462),
            data_re_in(15) => mul_re_out(463),
            data_re_in(16) => mul_re_out(464),
            data_re_in(17) => mul_re_out(465),
            data_re_in(18) => mul_re_out(466),
            data_re_in(19) => mul_re_out(467),
            data_re_in(20) => mul_re_out(468),
            data_re_in(21) => mul_re_out(469),
            data_re_in(22) => mul_re_out(470),
            data_re_in(23) => mul_re_out(471),
            data_re_in(24) => mul_re_out(472),
            data_re_in(25) => mul_re_out(473),
            data_re_in(26) => mul_re_out(474),
            data_re_in(27) => mul_re_out(475),
            data_re_in(28) => mul_re_out(476),
            data_re_in(29) => mul_re_out(477),
            data_re_in(30) => mul_re_out(478),
            data_re_in(31) => mul_re_out(479),
            data_im_in(0) => mul_im_out(448),
            data_im_in(1) => mul_im_out(449),
            data_im_in(2) => mul_im_out(450),
            data_im_in(3) => mul_im_out(451),
            data_im_in(4) => mul_im_out(452),
            data_im_in(5) => mul_im_out(453),
            data_im_in(6) => mul_im_out(454),
            data_im_in(7) => mul_im_out(455),
            data_im_in(8) => mul_im_out(456),
            data_im_in(9) => mul_im_out(457),
            data_im_in(10) => mul_im_out(458),
            data_im_in(11) => mul_im_out(459),
            data_im_in(12) => mul_im_out(460),
            data_im_in(13) => mul_im_out(461),
            data_im_in(14) => mul_im_out(462),
            data_im_in(15) => mul_im_out(463),
            data_im_in(16) => mul_im_out(464),
            data_im_in(17) => mul_im_out(465),
            data_im_in(18) => mul_im_out(466),
            data_im_in(19) => mul_im_out(467),
            data_im_in(20) => mul_im_out(468),
            data_im_in(21) => mul_im_out(469),
            data_im_in(22) => mul_im_out(470),
            data_im_in(23) => mul_im_out(471),
            data_im_in(24) => mul_im_out(472),
            data_im_in(25) => mul_im_out(473),
            data_im_in(26) => mul_im_out(474),
            data_im_in(27) => mul_im_out(475),
            data_im_in(28) => mul_im_out(476),
            data_im_in(29) => mul_im_out(477),
            data_im_in(30) => mul_im_out(478),
            data_im_in(31) => mul_im_out(479),
            data_re_out(0) => data_re_out(14),
            data_re_out(1) => data_re_out(30),
            data_re_out(2) => data_re_out(46),
            data_re_out(3) => data_re_out(62),
            data_re_out(4) => data_re_out(78),
            data_re_out(5) => data_re_out(94),
            data_re_out(6) => data_re_out(110),
            data_re_out(7) => data_re_out(126),
            data_re_out(8) => data_re_out(142),
            data_re_out(9) => data_re_out(158),
            data_re_out(10) => data_re_out(174),
            data_re_out(11) => data_re_out(190),
            data_re_out(12) => data_re_out(206),
            data_re_out(13) => data_re_out(222),
            data_re_out(14) => data_re_out(238),
            data_re_out(15) => data_re_out(254),
            data_re_out(16) => data_re_out(270),
            data_re_out(17) => data_re_out(286),
            data_re_out(18) => data_re_out(302),
            data_re_out(19) => data_re_out(318),
            data_re_out(20) => data_re_out(334),
            data_re_out(21) => data_re_out(350),
            data_re_out(22) => data_re_out(366),
            data_re_out(23) => data_re_out(382),
            data_re_out(24) => data_re_out(398),
            data_re_out(25) => data_re_out(414),
            data_re_out(26) => data_re_out(430),
            data_re_out(27) => data_re_out(446),
            data_re_out(28) => data_re_out(462),
            data_re_out(29) => data_re_out(478),
            data_re_out(30) => data_re_out(494),
            data_re_out(31) => data_re_out(510),
            data_im_out(0) => data_im_out(14),
            data_im_out(1) => data_im_out(30),
            data_im_out(2) => data_im_out(46),
            data_im_out(3) => data_im_out(62),
            data_im_out(4) => data_im_out(78),
            data_im_out(5) => data_im_out(94),
            data_im_out(6) => data_im_out(110),
            data_im_out(7) => data_im_out(126),
            data_im_out(8) => data_im_out(142),
            data_im_out(9) => data_im_out(158),
            data_im_out(10) => data_im_out(174),
            data_im_out(11) => data_im_out(190),
            data_im_out(12) => data_im_out(206),
            data_im_out(13) => data_im_out(222),
            data_im_out(14) => data_im_out(238),
            data_im_out(15) => data_im_out(254),
            data_im_out(16) => data_im_out(270),
            data_im_out(17) => data_im_out(286),
            data_im_out(18) => data_im_out(302),
            data_im_out(19) => data_im_out(318),
            data_im_out(20) => data_im_out(334),
            data_im_out(21) => data_im_out(350),
            data_im_out(22) => data_im_out(366),
            data_im_out(23) => data_im_out(382),
            data_im_out(24) => data_im_out(398),
            data_im_out(25) => data_im_out(414),
            data_im_out(26) => data_im_out(430),
            data_im_out(27) => data_im_out(446),
            data_im_out(28) => data_im_out(462),
            data_im_out(29) => data_im_out(478),
            data_im_out(30) => data_im_out(494),
            data_im_out(31) => data_im_out(510)
        );           

    URFFT_PT32_15 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(480),
            data_re_in(1) => mul_re_out(481),
            data_re_in(2) => mul_re_out(482),
            data_re_in(3) => mul_re_out(483),
            data_re_in(4) => mul_re_out(484),
            data_re_in(5) => mul_re_out(485),
            data_re_in(6) => mul_re_out(486),
            data_re_in(7) => mul_re_out(487),
            data_re_in(8) => mul_re_out(488),
            data_re_in(9) => mul_re_out(489),
            data_re_in(10) => mul_re_out(490),
            data_re_in(11) => mul_re_out(491),
            data_re_in(12) => mul_re_out(492),
            data_re_in(13) => mul_re_out(493),
            data_re_in(14) => mul_re_out(494),
            data_re_in(15) => mul_re_out(495),
            data_re_in(16) => mul_re_out(496),
            data_re_in(17) => mul_re_out(497),
            data_re_in(18) => mul_re_out(498),
            data_re_in(19) => mul_re_out(499),
            data_re_in(20) => mul_re_out(500),
            data_re_in(21) => mul_re_out(501),
            data_re_in(22) => mul_re_out(502),
            data_re_in(23) => mul_re_out(503),
            data_re_in(24) => mul_re_out(504),
            data_re_in(25) => mul_re_out(505),
            data_re_in(26) => mul_re_out(506),
            data_re_in(27) => mul_re_out(507),
            data_re_in(28) => mul_re_out(508),
            data_re_in(29) => mul_re_out(509),
            data_re_in(30) => mul_re_out(510),
            data_re_in(31) => mul_re_out(511),
            data_im_in(0) => mul_im_out(480),
            data_im_in(1) => mul_im_out(481),
            data_im_in(2) => mul_im_out(482),
            data_im_in(3) => mul_im_out(483),
            data_im_in(4) => mul_im_out(484),
            data_im_in(5) => mul_im_out(485),
            data_im_in(6) => mul_im_out(486),
            data_im_in(7) => mul_im_out(487),
            data_im_in(8) => mul_im_out(488),
            data_im_in(9) => mul_im_out(489),
            data_im_in(10) => mul_im_out(490),
            data_im_in(11) => mul_im_out(491),
            data_im_in(12) => mul_im_out(492),
            data_im_in(13) => mul_im_out(493),
            data_im_in(14) => mul_im_out(494),
            data_im_in(15) => mul_im_out(495),
            data_im_in(16) => mul_im_out(496),
            data_im_in(17) => mul_im_out(497),
            data_im_in(18) => mul_im_out(498),
            data_im_in(19) => mul_im_out(499),
            data_im_in(20) => mul_im_out(500),
            data_im_in(21) => mul_im_out(501),
            data_im_in(22) => mul_im_out(502),
            data_im_in(23) => mul_im_out(503),
            data_im_in(24) => mul_im_out(504),
            data_im_in(25) => mul_im_out(505),
            data_im_in(26) => mul_im_out(506),
            data_im_in(27) => mul_im_out(507),
            data_im_in(28) => mul_im_out(508),
            data_im_in(29) => mul_im_out(509),
            data_im_in(30) => mul_im_out(510),
            data_im_in(31) => mul_im_out(511),
            data_re_out(0) => data_re_out(15),
            data_re_out(1) => data_re_out(31),
            data_re_out(2) => data_re_out(47),
            data_re_out(3) => data_re_out(63),
            data_re_out(4) => data_re_out(79),
            data_re_out(5) => data_re_out(95),
            data_re_out(6) => data_re_out(111),
            data_re_out(7) => data_re_out(127),
            data_re_out(8) => data_re_out(143),
            data_re_out(9) => data_re_out(159),
            data_re_out(10) => data_re_out(175),
            data_re_out(11) => data_re_out(191),
            data_re_out(12) => data_re_out(207),
            data_re_out(13) => data_re_out(223),
            data_re_out(14) => data_re_out(239),
            data_re_out(15) => data_re_out(255),
            data_re_out(16) => data_re_out(271),
            data_re_out(17) => data_re_out(287),
            data_re_out(18) => data_re_out(303),
            data_re_out(19) => data_re_out(319),
            data_re_out(20) => data_re_out(335),
            data_re_out(21) => data_re_out(351),
            data_re_out(22) => data_re_out(367),
            data_re_out(23) => data_re_out(383),
            data_re_out(24) => data_re_out(399),
            data_re_out(25) => data_re_out(415),
            data_re_out(26) => data_re_out(431),
            data_re_out(27) => data_re_out(447),
            data_re_out(28) => data_re_out(463),
            data_re_out(29) => data_re_out(479),
            data_re_out(30) => data_re_out(495),
            data_re_out(31) => data_re_out(511),
            data_im_out(0) => data_im_out(15),
            data_im_out(1) => data_im_out(31),
            data_im_out(2) => data_im_out(47),
            data_im_out(3) => data_im_out(63),
            data_im_out(4) => data_im_out(79),
            data_im_out(5) => data_im_out(95),
            data_im_out(6) => data_im_out(111),
            data_im_out(7) => data_im_out(127),
            data_im_out(8) => data_im_out(143),
            data_im_out(9) => data_im_out(159),
            data_im_out(10) => data_im_out(175),
            data_im_out(11) => data_im_out(191),
            data_im_out(12) => data_im_out(207),
            data_im_out(13) => data_im_out(223),
            data_im_out(14) => data_im_out(239),
            data_im_out(15) => data_im_out(255),
            data_im_out(16) => data_im_out(271),
            data_im_out(17) => data_im_out(287),
            data_im_out(18) => data_im_out(303),
            data_im_out(19) => data_im_out(319),
            data_im_out(20) => data_im_out(335),
            data_im_out(21) => data_im_out(351),
            data_im_out(22) => data_im_out(367),
            data_im_out(23) => data_im_out(383),
            data_im_out(24) => data_im_out(399),
            data_im_out(25) => data_im_out(415),
            data_im_out(26) => data_im_out(431),
            data_im_out(27) => data_im_out(447),
            data_im_out(28) => data_im_out(463),
            data_im_out(29) => data_im_out(479),
            data_im_out(30) => data_im_out(495),
            data_im_out(31) => data_im_out(511)
        );           


    --- multipliers
 
    UMUL_0 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(0),
            data_im_in => first_stage_im_out(0),
            data_re_out => mul_re_out(0),
            data_im_out => mul_im_out(0)
        );

 
    UMUL_1 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1),
            data_im_in => first_stage_im_out(1),
            data_re_out => mul_re_out(1),
            data_im_out => mul_im_out(1)
        );

 
    UMUL_2 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2),
            data_im_in => first_stage_im_out(2),
            data_re_out => mul_re_out(2),
            data_im_out => mul_im_out(2)
        );

 
    UMUL_3 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(3),
            data_im_in => first_stage_im_out(3),
            data_re_out => mul_re_out(3),
            data_im_out => mul_im_out(3)
        );

 
    UMUL_4 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(4),
            data_im_in => first_stage_im_out(4),
            data_re_out => mul_re_out(4),
            data_im_out => mul_im_out(4)
        );

 
    UMUL_5 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(5),
            data_im_in => first_stage_im_out(5),
            data_re_out => mul_re_out(5),
            data_im_out => mul_im_out(5)
        );

 
    UMUL_6 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(6),
            data_im_in => first_stage_im_out(6),
            data_re_out => mul_re_out(6),
            data_im_out => mul_im_out(6)
        );

 
    UMUL_7 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(7),
            data_im_in => first_stage_im_out(7),
            data_re_out => mul_re_out(7),
            data_im_out => mul_im_out(7)
        );

 
    UMUL_8 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(8),
            data_im_in => first_stage_im_out(8),
            data_re_out => mul_re_out(8),
            data_im_out => mul_im_out(8)
        );

 
    UMUL_9 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(9),
            data_im_in => first_stage_im_out(9),
            data_re_out => mul_re_out(9),
            data_im_out => mul_im_out(9)
        );

 
    UMUL_10 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(10),
            data_im_in => first_stage_im_out(10),
            data_re_out => mul_re_out(10),
            data_im_out => mul_im_out(10)
        );

 
    UMUL_11 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(11),
            data_im_in => first_stage_im_out(11),
            data_re_out => mul_re_out(11),
            data_im_out => mul_im_out(11)
        );

 
    UMUL_12 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(12),
            data_im_in => first_stage_im_out(12),
            data_re_out => mul_re_out(12),
            data_im_out => mul_im_out(12)
        );

 
    UMUL_13 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(13),
            data_im_in => first_stage_im_out(13),
            data_re_out => mul_re_out(13),
            data_im_out => mul_im_out(13)
        );

 
    UMUL_14 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(14),
            data_im_in => first_stage_im_out(14),
            data_re_out => mul_re_out(14),
            data_im_out => mul_im_out(14)
        );

 
    UMUL_15 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(15),
            data_im_in => first_stage_im_out(15),
            data_re_out => mul_re_out(15),
            data_im_out => mul_im_out(15)
        );

 
    UMUL_16 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(16),
            data_im_in => first_stage_im_out(16),
            data_re_out => mul_re_out(16),
            data_im_out => mul_im_out(16)
        );

 
    UMUL_17 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(17),
            data_im_in => first_stage_im_out(17),
            data_re_out => mul_re_out(17),
            data_im_out => mul_im_out(17)
        );

 
    UMUL_18 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(18),
            data_im_in => first_stage_im_out(18),
            data_re_out => mul_re_out(18),
            data_im_out => mul_im_out(18)
        );

 
    UMUL_19 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(19),
            data_im_in => first_stage_im_out(19),
            data_re_out => mul_re_out(19),
            data_im_out => mul_im_out(19)
        );

 
    UMUL_20 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(20),
            data_im_in => first_stage_im_out(20),
            data_re_out => mul_re_out(20),
            data_im_out => mul_im_out(20)
        );

 
    UMUL_21 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(21),
            data_im_in => first_stage_im_out(21),
            data_re_out => mul_re_out(21),
            data_im_out => mul_im_out(21)
        );

 
    UMUL_22 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(22),
            data_im_in => first_stage_im_out(22),
            data_re_out => mul_re_out(22),
            data_im_out => mul_im_out(22)
        );

 
    UMUL_23 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(23),
            data_im_in => first_stage_im_out(23),
            data_re_out => mul_re_out(23),
            data_im_out => mul_im_out(23)
        );

 
    UMUL_24 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(24),
            data_im_in => first_stage_im_out(24),
            data_re_out => mul_re_out(24),
            data_im_out => mul_im_out(24)
        );

 
    UMUL_25 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(25),
            data_im_in => first_stage_im_out(25),
            data_re_out => mul_re_out(25),
            data_im_out => mul_im_out(25)
        );

 
    UMUL_26 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(26),
            data_im_in => first_stage_im_out(26),
            data_re_out => mul_re_out(26),
            data_im_out => mul_im_out(26)
        );

 
    UMUL_27 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(27),
            data_im_in => first_stage_im_out(27),
            data_re_out => mul_re_out(27),
            data_im_out => mul_im_out(27)
        );

 
    UMUL_28 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(28),
            data_im_in => first_stage_im_out(28),
            data_re_out => mul_re_out(28),
            data_im_out => mul_im_out(28)
        );

 
    UMUL_29 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(29),
            data_im_in => first_stage_im_out(29),
            data_re_out => mul_re_out(29),
            data_im_out => mul_im_out(29)
        );

 
    UMUL_30 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(30),
            data_im_in => first_stage_im_out(30),
            data_re_out => mul_re_out(30),
            data_im_out => mul_im_out(30)
        );

 
    UMUL_31 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(31),
            data_im_in => first_stage_im_out(31),
            data_re_out => mul_re_out(31),
            data_im_out => mul_im_out(31)
        );

 
    UMUL_32 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(32),
            data_im_in => first_stage_im_out(32),
            data_re_out => mul_re_out(32),
            data_im_out => mul_im_out(32)
        );

 
    UMUL_33 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(33),
            data_im_in => first_stage_im_out(33),
            re_multiplicator => re_multiplicator(33), ---  0.999938964844
            im_multiplicator => im_multiplicator(33), --- j-0.0122680664062
            data_re_out => mul_re_out(33),
            data_im_out => mul_im_out(33)
        );

 
    UMUL_34 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(34),
            data_im_in => first_stage_im_out(34),
            re_multiplicator => re_multiplicator(34), ---  0.999694824219
            im_multiplicator => im_multiplicator(34), --- j-0.0245361328125
            data_re_out => mul_re_out(34),
            data_im_out => mul_im_out(34)
        );

 
    UMUL_35 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(35),
            data_im_in => first_stage_im_out(35),
            re_multiplicator => re_multiplicator(35), ---  0.999328613281
            im_multiplicator => im_multiplicator(35), --- j-0.0368041992188
            data_re_out => mul_re_out(35),
            data_im_out => mul_im_out(35)
        );

 
    UMUL_36 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(36),
            data_im_in => first_stage_im_out(36),
            re_multiplicator => re_multiplicator(36), ---  0.998779296875
            im_multiplicator => im_multiplicator(36), --- j-0.049072265625
            data_re_out => mul_re_out(36),
            data_im_out => mul_im_out(36)
        );

 
    UMUL_37 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(37),
            data_im_in => first_stage_im_out(37),
            re_multiplicator => re_multiplicator(37), ---  0.998107910156
            im_multiplicator => im_multiplicator(37), --- j-0.0613403320312
            data_re_out => mul_re_out(37),
            data_im_out => mul_im_out(37)
        );

 
    UMUL_38 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(38),
            data_im_in => first_stage_im_out(38),
            re_multiplicator => re_multiplicator(38), ---  0.997314453125
            im_multiplicator => im_multiplicator(38), --- j-0.0735473632812
            data_re_out => mul_re_out(38),
            data_im_out => mul_im_out(38)
        );

 
    UMUL_39 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(39),
            data_im_in => first_stage_im_out(39),
            re_multiplicator => re_multiplicator(39), ---  0.996337890625
            im_multiplicator => im_multiplicator(39), --- j-0.0858154296875
            data_re_out => mul_re_out(39),
            data_im_out => mul_im_out(39)
        );

 
    UMUL_40 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(40),
            data_im_in => first_stage_im_out(40),
            re_multiplicator => re_multiplicator(40), ---  0.995178222656
            im_multiplicator => im_multiplicator(40), --- j-0.0980224609375
            data_re_out => mul_re_out(40),
            data_im_out => mul_im_out(40)
        );

 
    UMUL_41 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(41),
            data_im_in => first_stage_im_out(41),
            re_multiplicator => re_multiplicator(41), ---  0.993896484375
            im_multiplicator => im_multiplicator(41), --- j-0.110229492188
            data_re_out => mul_re_out(41),
            data_im_out => mul_im_out(41)
        );

 
    UMUL_42 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(42),
            data_im_in => first_stage_im_out(42),
            re_multiplicator => re_multiplicator(42), ---  0.992492675781
            im_multiplicator => im_multiplicator(42), --- j-0.122436523438
            data_re_out => mul_re_out(42),
            data_im_out => mul_im_out(42)
        );

 
    UMUL_43 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(43),
            data_im_in => first_stage_im_out(43),
            re_multiplicator => re_multiplicator(43), ---  0.990905761719
            im_multiplicator => im_multiplicator(43), --- j-0.134582519531
            data_re_out => mul_re_out(43),
            data_im_out => mul_im_out(43)
        );

 
    UMUL_44 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(44),
            data_im_in => first_stage_im_out(44),
            re_multiplicator => re_multiplicator(44), ---  0.989196777344
            im_multiplicator => im_multiplicator(44), --- j-0.146728515625
            data_re_out => mul_re_out(44),
            data_im_out => mul_im_out(44)
        );

 
    UMUL_45 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(45),
            data_im_in => first_stage_im_out(45),
            re_multiplicator => re_multiplicator(45), ---  0.9873046875
            im_multiplicator => im_multiplicator(45), --- j-0.158874511719
            data_re_out => mul_re_out(45),
            data_im_out => mul_im_out(45)
        );

 
    UMUL_46 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(46),
            data_im_in => first_stage_im_out(46),
            re_multiplicator => re_multiplicator(46), ---  0.985290527344
            im_multiplicator => im_multiplicator(46), --- j-0.170959472656
            data_re_out => mul_re_out(46),
            data_im_out => mul_im_out(46)
        );

 
    UMUL_47 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(47),
            data_im_in => first_stage_im_out(47),
            re_multiplicator => re_multiplicator(47), ---  0.983093261719
            im_multiplicator => im_multiplicator(47), --- j-0.183044433594
            data_re_out => mul_re_out(47),
            data_im_out => mul_im_out(47)
        );

 
    UMUL_48 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(48),
            data_im_in => first_stage_im_out(48),
            re_multiplicator => re_multiplicator(48), ---  0.980773925781
            im_multiplicator => im_multiplicator(48), --- j-0.195068359375
            data_re_out => mul_re_out(48),
            data_im_out => mul_im_out(48)
        );

 
    UMUL_49 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(49),
            data_im_in => first_stage_im_out(49),
            re_multiplicator => re_multiplicator(49), ---  0.978332519531
            im_multiplicator => im_multiplicator(49), --- j-0.207092285156
            data_re_out => mul_re_out(49),
            data_im_out => mul_im_out(49)
        );

 
    UMUL_50 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(50),
            data_im_in => first_stage_im_out(50),
            re_multiplicator => re_multiplicator(50), ---  0.975708007812
            im_multiplicator => im_multiplicator(50), --- j-0.219116210938
            data_re_out => mul_re_out(50),
            data_im_out => mul_im_out(50)
        );

 
    UMUL_51 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(51),
            data_im_in => first_stage_im_out(51),
            re_multiplicator => re_multiplicator(51), ---  0.972961425781
            im_multiplicator => im_multiplicator(51), --- j-0.231079101562
            data_re_out => mul_re_out(51),
            data_im_out => mul_im_out(51)
        );

 
    UMUL_52 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(52),
            data_im_in => first_stage_im_out(52),
            re_multiplicator => re_multiplicator(52), ---  0.970031738281
            im_multiplicator => im_multiplicator(52), --- j-0.242980957031
            data_re_out => mul_re_out(52),
            data_im_out => mul_im_out(52)
        );

 
    UMUL_53 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(53),
            data_im_in => first_stage_im_out(53),
            re_multiplicator => re_multiplicator(53), ---  0.966979980469
            im_multiplicator => im_multiplicator(53), --- j-0.2548828125
            data_re_out => mul_re_out(53),
            data_im_out => mul_im_out(53)
        );

 
    UMUL_54 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(54),
            data_im_in => first_stage_im_out(54),
            re_multiplicator => re_multiplicator(54), ---  0.963806152344
            im_multiplicator => im_multiplicator(54), --- j-0.266723632812
            data_re_out => mul_re_out(54),
            data_im_out => mul_im_out(54)
        );

 
    UMUL_55 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(55),
            data_im_in => first_stage_im_out(55),
            re_multiplicator => re_multiplicator(55), ---  0.96044921875
            im_multiplicator => im_multiplicator(55), --- j-0.278503417969
            data_re_out => mul_re_out(55),
            data_im_out => mul_im_out(55)
        );

 
    UMUL_56 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(56),
            data_im_in => first_stage_im_out(56),
            re_multiplicator => re_multiplicator(56), ---  0.956970214844
            im_multiplicator => im_multiplicator(56), --- j-0.290283203125
            data_re_out => mul_re_out(56),
            data_im_out => mul_im_out(56)
        );

 
    UMUL_57 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(57),
            data_im_in => first_stage_im_out(57),
            re_multiplicator => re_multiplicator(57), ---  0.953308105469
            im_multiplicator => im_multiplicator(57), --- j-0.302001953125
            data_re_out => mul_re_out(57),
            data_im_out => mul_im_out(57)
        );

 
    UMUL_58 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(58),
            data_im_in => first_stage_im_out(58),
            re_multiplicator => re_multiplicator(58), ---  0.949523925781
            im_multiplicator => im_multiplicator(58), --- j-0.313659667969
            data_re_out => mul_re_out(58),
            data_im_out => mul_im_out(58)
        );

 
    UMUL_59 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(59),
            data_im_in => first_stage_im_out(59),
            re_multiplicator => re_multiplicator(59), ---  0.945617675781
            im_multiplicator => im_multiplicator(59), --- j-0.325317382812
            data_re_out => mul_re_out(59),
            data_im_out => mul_im_out(59)
        );

 
    UMUL_60 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(60),
            data_im_in => first_stage_im_out(60),
            re_multiplicator => re_multiplicator(60), ---  0.941528320312
            im_multiplicator => im_multiplicator(60), --- j-0.3369140625
            data_re_out => mul_re_out(60),
            data_im_out => mul_im_out(60)
        );

 
    UMUL_61 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(61),
            data_im_in => first_stage_im_out(61),
            re_multiplicator => re_multiplicator(61), ---  0.937316894531
            im_multiplicator => im_multiplicator(61), --- j-0.348388671875
            data_re_out => mul_re_out(61),
            data_im_out => mul_im_out(61)
        );

 
    UMUL_62 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(62),
            data_im_in => first_stage_im_out(62),
            re_multiplicator => re_multiplicator(62), ---  0.932983398438
            im_multiplicator => im_multiplicator(62), --- j-0.359924316406
            data_re_out => mul_re_out(62),
            data_im_out => mul_im_out(62)
        );

 
    UMUL_63 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(63),
            data_im_in => first_stage_im_out(63),
            re_multiplicator => re_multiplicator(63), ---  0.928527832031
            im_multiplicator => im_multiplicator(63), --- j-0.371337890625
            data_re_out => mul_re_out(63),
            data_im_out => mul_im_out(63)
        );

 
    UMUL_64 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(64),
            data_im_in => first_stage_im_out(64),
            data_re_out => mul_re_out(64),
            data_im_out => mul_im_out(64)
        );

 
    UMUL_65 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(65),
            data_im_in => first_stage_im_out(65),
            re_multiplicator => re_multiplicator(65), ---  0.999694824219
            im_multiplicator => im_multiplicator(65), --- j-0.0245361328125
            data_re_out => mul_re_out(65),
            data_im_out => mul_im_out(65)
        );

 
    UMUL_66 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(66),
            data_im_in => first_stage_im_out(66),
            re_multiplicator => re_multiplicator(66), ---  0.998779296875
            im_multiplicator => im_multiplicator(66), --- j-0.049072265625
            data_re_out => mul_re_out(66),
            data_im_out => mul_im_out(66)
        );

 
    UMUL_67 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(67),
            data_im_in => first_stage_im_out(67),
            re_multiplicator => re_multiplicator(67), ---  0.997314453125
            im_multiplicator => im_multiplicator(67), --- j-0.0735473632812
            data_re_out => mul_re_out(67),
            data_im_out => mul_im_out(67)
        );

 
    UMUL_68 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(68),
            data_im_in => first_stage_im_out(68),
            re_multiplicator => re_multiplicator(68), ---  0.995178222656
            im_multiplicator => im_multiplicator(68), --- j-0.0980224609375
            data_re_out => mul_re_out(68),
            data_im_out => mul_im_out(68)
        );

 
    UMUL_69 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(69),
            data_im_in => first_stage_im_out(69),
            re_multiplicator => re_multiplicator(69), ---  0.992492675781
            im_multiplicator => im_multiplicator(69), --- j-0.122436523438
            data_re_out => mul_re_out(69),
            data_im_out => mul_im_out(69)
        );

 
    UMUL_70 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(70),
            data_im_in => first_stage_im_out(70),
            re_multiplicator => re_multiplicator(70), ---  0.989196777344
            im_multiplicator => im_multiplicator(70), --- j-0.146728515625
            data_re_out => mul_re_out(70),
            data_im_out => mul_im_out(70)
        );

 
    UMUL_71 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(71),
            data_im_in => first_stage_im_out(71),
            re_multiplicator => re_multiplicator(71), ---  0.985290527344
            im_multiplicator => im_multiplicator(71), --- j-0.170959472656
            data_re_out => mul_re_out(71),
            data_im_out => mul_im_out(71)
        );

 
    UMUL_72 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(72),
            data_im_in => first_stage_im_out(72),
            re_multiplicator => re_multiplicator(72), ---  0.980773925781
            im_multiplicator => im_multiplicator(72), --- j-0.195068359375
            data_re_out => mul_re_out(72),
            data_im_out => mul_im_out(72)
        );

 
    UMUL_73 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(73),
            data_im_in => first_stage_im_out(73),
            re_multiplicator => re_multiplicator(73), ---  0.975708007812
            im_multiplicator => im_multiplicator(73), --- j-0.219116210938
            data_re_out => mul_re_out(73),
            data_im_out => mul_im_out(73)
        );

 
    UMUL_74 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(74),
            data_im_in => first_stage_im_out(74),
            re_multiplicator => re_multiplicator(74), ---  0.970031738281
            im_multiplicator => im_multiplicator(74), --- j-0.242980957031
            data_re_out => mul_re_out(74),
            data_im_out => mul_im_out(74)
        );

 
    UMUL_75 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(75),
            data_im_in => first_stage_im_out(75),
            re_multiplicator => re_multiplicator(75), ---  0.963806152344
            im_multiplicator => im_multiplicator(75), --- j-0.266723632812
            data_re_out => mul_re_out(75),
            data_im_out => mul_im_out(75)
        );

 
    UMUL_76 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(76),
            data_im_in => first_stage_im_out(76),
            re_multiplicator => re_multiplicator(76), ---  0.956970214844
            im_multiplicator => im_multiplicator(76), --- j-0.290283203125
            data_re_out => mul_re_out(76),
            data_im_out => mul_im_out(76)
        );

 
    UMUL_77 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(77),
            data_im_in => first_stage_im_out(77),
            re_multiplicator => re_multiplicator(77), ---  0.949523925781
            im_multiplicator => im_multiplicator(77), --- j-0.313659667969
            data_re_out => mul_re_out(77),
            data_im_out => mul_im_out(77)
        );

 
    UMUL_78 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(78),
            data_im_in => first_stage_im_out(78),
            re_multiplicator => re_multiplicator(78), ---  0.941528320312
            im_multiplicator => im_multiplicator(78), --- j-0.3369140625
            data_re_out => mul_re_out(78),
            data_im_out => mul_im_out(78)
        );

 
    UMUL_79 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(79),
            data_im_in => first_stage_im_out(79),
            re_multiplicator => re_multiplicator(79), ---  0.932983398438
            im_multiplicator => im_multiplicator(79), --- j-0.359924316406
            data_re_out => mul_re_out(79),
            data_im_out => mul_im_out(79)
        );

 
    UMUL_80 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(80),
            data_im_in => first_stage_im_out(80),
            re_multiplicator => re_multiplicator(80), ---  0.923889160156
            im_multiplicator => im_multiplicator(80), --- j-0.382690429688
            data_re_out => mul_re_out(80),
            data_im_out => mul_im_out(80)
        );

 
    UMUL_81 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(81),
            data_im_in => first_stage_im_out(81),
            re_multiplicator => re_multiplicator(81), ---  0.914184570312
            im_multiplicator => im_multiplicator(81), --- j-0.405212402344
            data_re_out => mul_re_out(81),
            data_im_out => mul_im_out(81)
        );

 
    UMUL_82 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(82),
            data_im_in => first_stage_im_out(82),
            re_multiplicator => re_multiplicator(82), ---  0.903991699219
            im_multiplicator => im_multiplicator(82), --- j-0.427551269531
            data_re_out => mul_re_out(82),
            data_im_out => mul_im_out(82)
        );

 
    UMUL_83 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(83),
            data_im_in => first_stage_im_out(83),
            re_multiplicator => re_multiplicator(83), ---  0.893249511719
            im_multiplicator => im_multiplicator(83), --- j-0.449584960938
            data_re_out => mul_re_out(83),
            data_im_out => mul_im_out(83)
        );

 
    UMUL_84 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(84),
            data_im_in => first_stage_im_out(84),
            re_multiplicator => re_multiplicator(84), ---  0.881896972656
            im_multiplicator => im_multiplicator(84), --- j-0.471374511719
            data_re_out => mul_re_out(84),
            data_im_out => mul_im_out(84)
        );

 
    UMUL_85 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(85),
            data_im_in => first_stage_im_out(85),
            re_multiplicator => re_multiplicator(85), ---  0.8701171875
            im_multiplicator => im_multiplicator(85), --- j-0.492919921875
            data_re_out => mul_re_out(85),
            data_im_out => mul_im_out(85)
        );

 
    UMUL_86 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(86),
            data_im_in => first_stage_im_out(86),
            re_multiplicator => re_multiplicator(86), ---  0.857727050781
            im_multiplicator => im_multiplicator(86), --- j-0.514099121094
            data_re_out => mul_re_out(86),
            data_im_out => mul_im_out(86)
        );

 
    UMUL_87 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(87),
            data_im_in => first_stage_im_out(87),
            re_multiplicator => re_multiplicator(87), ---  0.844848632812
            im_multiplicator => im_multiplicator(87), --- j-0.534973144531
            data_re_out => mul_re_out(87),
            data_im_out => mul_im_out(87)
        );

 
    UMUL_88 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(88),
            data_im_in => first_stage_im_out(88),
            re_multiplicator => re_multiplicator(88), ---  0.831481933594
            im_multiplicator => im_multiplicator(88), --- j-0.555541992188
            data_re_out => mul_re_out(88),
            data_im_out => mul_im_out(88)
        );

 
    UMUL_89 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(89),
            data_im_in => first_stage_im_out(89),
            re_multiplicator => re_multiplicator(89), ---  0.817565917969
            im_multiplicator => im_multiplicator(89), --- j-0.575805664062
            data_re_out => mul_re_out(89),
            data_im_out => mul_im_out(89)
        );

 
    UMUL_90 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(90),
            data_im_in => first_stage_im_out(90),
            re_multiplicator => re_multiplicator(90), ---  0.80322265625
            im_multiplicator => im_multiplicator(90), --- j-0.595703125
            data_re_out => mul_re_out(90),
            data_im_out => mul_im_out(90)
        );

 
    UMUL_91 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(91),
            data_im_in => first_stage_im_out(91),
            re_multiplicator => re_multiplicator(91), ---  0.788330078125
            im_multiplicator => im_multiplicator(91), --- j-0.615234375
            data_re_out => mul_re_out(91),
            data_im_out => mul_im_out(91)
        );

 
    UMUL_92 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(92),
            data_im_in => first_stage_im_out(92),
            re_multiplicator => re_multiplicator(92), ---  0.773010253906
            im_multiplicator => im_multiplicator(92), --- j-0.634399414062
            data_re_out => mul_re_out(92),
            data_im_out => mul_im_out(92)
        );

 
    UMUL_93 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(93),
            data_im_in => first_stage_im_out(93),
            re_multiplicator => re_multiplicator(93), ---  0.757202148438
            im_multiplicator => im_multiplicator(93), --- j-0.653198242188
            data_re_out => mul_re_out(93),
            data_im_out => mul_im_out(93)
        );

 
    UMUL_94 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(94),
            data_im_in => first_stage_im_out(94),
            re_multiplicator => re_multiplicator(94), ---  0.740966796875
            im_multiplicator => im_multiplicator(94), --- j-0.671569824219
            data_re_out => mul_re_out(94),
            data_im_out => mul_im_out(94)
        );

 
    UMUL_95 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(95),
            data_im_in => first_stage_im_out(95),
            re_multiplicator => re_multiplicator(95), ---  0.724243164062
            im_multiplicator => im_multiplicator(95), --- j-0.689514160156
            data_re_out => mul_re_out(95),
            data_im_out => mul_im_out(95)
        );

 
    UMUL_96 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(96),
            data_im_in => first_stage_im_out(96),
            data_re_out => mul_re_out(96),
            data_im_out => mul_im_out(96)
        );

 
    UMUL_97 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(97),
            data_im_in => first_stage_im_out(97),
            re_multiplicator => re_multiplicator(97), ---  0.999328613281
            im_multiplicator => im_multiplicator(97), --- j-0.0368041992188
            data_re_out => mul_re_out(97),
            data_im_out => mul_im_out(97)
        );

 
    UMUL_98 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(98),
            data_im_in => first_stage_im_out(98),
            re_multiplicator => re_multiplicator(98), ---  0.997314453125
            im_multiplicator => im_multiplicator(98), --- j-0.0735473632812
            data_re_out => mul_re_out(98),
            data_im_out => mul_im_out(98)
        );

 
    UMUL_99 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(99),
            data_im_in => first_stage_im_out(99),
            re_multiplicator => re_multiplicator(99), ---  0.993896484375
            im_multiplicator => im_multiplicator(99), --- j-0.110229492188
            data_re_out => mul_re_out(99),
            data_im_out => mul_im_out(99)
        );

 
    UMUL_100 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(100),
            data_im_in => first_stage_im_out(100),
            re_multiplicator => re_multiplicator(100), ---  0.989196777344
            im_multiplicator => im_multiplicator(100), --- j-0.146728515625
            data_re_out => mul_re_out(100),
            data_im_out => mul_im_out(100)
        );

 
    UMUL_101 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(101),
            data_im_in => first_stage_im_out(101),
            re_multiplicator => re_multiplicator(101), ---  0.983093261719
            im_multiplicator => im_multiplicator(101), --- j-0.183044433594
            data_re_out => mul_re_out(101),
            data_im_out => mul_im_out(101)
        );

 
    UMUL_102 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(102),
            data_im_in => first_stage_im_out(102),
            re_multiplicator => re_multiplicator(102), ---  0.975708007812
            im_multiplicator => im_multiplicator(102), --- j-0.219116210938
            data_re_out => mul_re_out(102),
            data_im_out => mul_im_out(102)
        );

 
    UMUL_103 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(103),
            data_im_in => first_stage_im_out(103),
            re_multiplicator => re_multiplicator(103), ---  0.966979980469
            im_multiplicator => im_multiplicator(103), --- j-0.2548828125
            data_re_out => mul_re_out(103),
            data_im_out => mul_im_out(103)
        );

 
    UMUL_104 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(104),
            data_im_in => first_stage_im_out(104),
            re_multiplicator => re_multiplicator(104), ---  0.956970214844
            im_multiplicator => im_multiplicator(104), --- j-0.290283203125
            data_re_out => mul_re_out(104),
            data_im_out => mul_im_out(104)
        );

 
    UMUL_105 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(105),
            data_im_in => first_stage_im_out(105),
            re_multiplicator => re_multiplicator(105), ---  0.945617675781
            im_multiplicator => im_multiplicator(105), --- j-0.325317382812
            data_re_out => mul_re_out(105),
            data_im_out => mul_im_out(105)
        );

 
    UMUL_106 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(106),
            data_im_in => first_stage_im_out(106),
            re_multiplicator => re_multiplicator(106), ---  0.932983398438
            im_multiplicator => im_multiplicator(106), --- j-0.359924316406
            data_re_out => mul_re_out(106),
            data_im_out => mul_im_out(106)
        );

 
    UMUL_107 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(107),
            data_im_in => first_stage_im_out(107),
            re_multiplicator => re_multiplicator(107), ---  0.919128417969
            im_multiplicator => im_multiplicator(107), --- j-0.393981933594
            data_re_out => mul_re_out(107),
            data_im_out => mul_im_out(107)
        );

 
    UMUL_108 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(108),
            data_im_in => first_stage_im_out(108),
            re_multiplicator => re_multiplicator(108), ---  0.903991699219
            im_multiplicator => im_multiplicator(108), --- j-0.427551269531
            data_re_out => mul_re_out(108),
            data_im_out => mul_im_out(108)
        );

 
    UMUL_109 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(109),
            data_im_in => first_stage_im_out(109),
            re_multiplicator => re_multiplicator(109), ---  0.887634277344
            im_multiplicator => im_multiplicator(109), --- j-0.460510253906
            data_re_out => mul_re_out(109),
            data_im_out => mul_im_out(109)
        );

 
    UMUL_110 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(110),
            data_im_in => first_stage_im_out(110),
            re_multiplicator => re_multiplicator(110), ---  0.8701171875
            im_multiplicator => im_multiplicator(110), --- j-0.492919921875
            data_re_out => mul_re_out(110),
            data_im_out => mul_im_out(110)
        );

 
    UMUL_111 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(111),
            data_im_in => first_stage_im_out(111),
            re_multiplicator => re_multiplicator(111), ---  0.851379394531
            im_multiplicator => im_multiplicator(111), --- j-0.524597167969
            data_re_out => mul_re_out(111),
            data_im_out => mul_im_out(111)
        );

 
    UMUL_112 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(112),
            data_im_in => first_stage_im_out(112),
            re_multiplicator => re_multiplicator(112), ---  0.831481933594
            im_multiplicator => im_multiplicator(112), --- j-0.555541992188
            data_re_out => mul_re_out(112),
            data_im_out => mul_im_out(112)
        );

 
    UMUL_113 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(113),
            data_im_in => first_stage_im_out(113),
            re_multiplicator => re_multiplicator(113), ---  0.810485839844
            im_multiplicator => im_multiplicator(113), --- j-0.585815429688
            data_re_out => mul_re_out(113),
            data_im_out => mul_im_out(113)
        );

 
    UMUL_114 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(114),
            data_im_in => first_stage_im_out(114),
            re_multiplicator => re_multiplicator(114), ---  0.788330078125
            im_multiplicator => im_multiplicator(114), --- j-0.615234375
            data_re_out => mul_re_out(114),
            data_im_out => mul_im_out(114)
        );

 
    UMUL_115 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(115),
            data_im_in => first_stage_im_out(115),
            re_multiplicator => re_multiplicator(115), ---  0.765197753906
            im_multiplicator => im_multiplicator(115), --- j-0.643859863281
            data_re_out => mul_re_out(115),
            data_im_out => mul_im_out(115)
        );

 
    UMUL_116 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(116),
            data_im_in => first_stage_im_out(116),
            re_multiplicator => re_multiplicator(116), ---  0.740966796875
            im_multiplicator => im_multiplicator(116), --- j-0.671569824219
            data_re_out => mul_re_out(116),
            data_im_out => mul_im_out(116)
        );

 
    UMUL_117 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(117),
            data_im_in => first_stage_im_out(117),
            re_multiplicator => re_multiplicator(117), ---  0.715759277344
            im_multiplicator => im_multiplicator(117), --- j-0.698364257812
            data_re_out => mul_re_out(117),
            data_im_out => mul_im_out(117)
        );

 
    UMUL_118 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(118),
            data_im_in => first_stage_im_out(118),
            re_multiplicator => re_multiplicator(118), ---  0.689514160156
            im_multiplicator => im_multiplicator(118), --- j-0.724243164062
            data_re_out => mul_re_out(118),
            data_im_out => mul_im_out(118)
        );

 
    UMUL_119 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(119),
            data_im_in => first_stage_im_out(119),
            re_multiplicator => re_multiplicator(119), ---  0.662414550781
            im_multiplicator => im_multiplicator(119), --- j-0.749145507812
            data_re_out => mul_re_out(119),
            data_im_out => mul_im_out(119)
        );

 
    UMUL_120 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(120),
            data_im_in => first_stage_im_out(120),
            re_multiplicator => re_multiplicator(120), ---  0.634399414062
            im_multiplicator => im_multiplicator(120), --- j-0.773010253906
            data_re_out => mul_re_out(120),
            data_im_out => mul_im_out(120)
        );

 
    UMUL_121 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(121),
            data_im_in => first_stage_im_out(121),
            re_multiplicator => re_multiplicator(121), ---  0.605529785156
            im_multiplicator => im_multiplicator(121), --- j-0.795837402344
            data_re_out => mul_re_out(121),
            data_im_out => mul_im_out(121)
        );

 
    UMUL_122 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(122),
            data_im_in => first_stage_im_out(122),
            re_multiplicator => re_multiplicator(122), ---  0.575805664062
            im_multiplicator => im_multiplicator(122), --- j-0.817565917969
            data_re_out => mul_re_out(122),
            data_im_out => mul_im_out(122)
        );

 
    UMUL_123 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(123),
            data_im_in => first_stage_im_out(123),
            re_multiplicator => re_multiplicator(123), ---  0.545349121094
            im_multiplicator => im_multiplicator(123), --- j-0.838195800781
            data_re_out => mul_re_out(123),
            data_im_out => mul_im_out(123)
        );

 
    UMUL_124 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(124),
            data_im_in => first_stage_im_out(124),
            re_multiplicator => re_multiplicator(124), ---  0.514099121094
            im_multiplicator => im_multiplicator(124), --- j-0.857727050781
            data_re_out => mul_re_out(124),
            data_im_out => mul_im_out(124)
        );

 
    UMUL_125 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(125),
            data_im_in => first_stage_im_out(125),
            re_multiplicator => re_multiplicator(125), ---  0.482177734375
            im_multiplicator => im_multiplicator(125), --- j-0.876098632812
            data_re_out => mul_re_out(125),
            data_im_out => mul_im_out(125)
        );

 
    UMUL_126 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(126),
            data_im_in => first_stage_im_out(126),
            re_multiplicator => re_multiplicator(126), ---  0.449584960938
            im_multiplicator => im_multiplicator(126), --- j-0.893249511719
            data_re_out => mul_re_out(126),
            data_im_out => mul_im_out(126)
        );

 
    UMUL_127 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(127),
            data_im_in => first_stage_im_out(127),
            re_multiplicator => re_multiplicator(127), ---  0.416442871094
            im_multiplicator => im_multiplicator(127), --- j-0.9091796875
            data_re_out => mul_re_out(127),
            data_im_out => mul_im_out(127)
        );

 
    UMUL_128 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(128),
            data_im_in => first_stage_im_out(128),
            data_re_out => mul_re_out(128),
            data_im_out => mul_im_out(128)
        );

 
    UMUL_129 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(129),
            data_im_in => first_stage_im_out(129),
            re_multiplicator => re_multiplicator(129), ---  0.998779296875
            im_multiplicator => im_multiplicator(129), --- j-0.049072265625
            data_re_out => mul_re_out(129),
            data_im_out => mul_im_out(129)
        );

 
    UMUL_130 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(130),
            data_im_in => first_stage_im_out(130),
            re_multiplicator => re_multiplicator(130), ---  0.995178222656
            im_multiplicator => im_multiplicator(130), --- j-0.0980224609375
            data_re_out => mul_re_out(130),
            data_im_out => mul_im_out(130)
        );

 
    UMUL_131 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(131),
            data_im_in => first_stage_im_out(131),
            re_multiplicator => re_multiplicator(131), ---  0.989196777344
            im_multiplicator => im_multiplicator(131), --- j-0.146728515625
            data_re_out => mul_re_out(131),
            data_im_out => mul_im_out(131)
        );

 
    UMUL_132 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(132),
            data_im_in => first_stage_im_out(132),
            re_multiplicator => re_multiplicator(132), ---  0.980773925781
            im_multiplicator => im_multiplicator(132), --- j-0.195068359375
            data_re_out => mul_re_out(132),
            data_im_out => mul_im_out(132)
        );

 
    UMUL_133 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(133),
            data_im_in => first_stage_im_out(133),
            re_multiplicator => re_multiplicator(133), ---  0.970031738281
            im_multiplicator => im_multiplicator(133), --- j-0.242980957031
            data_re_out => mul_re_out(133),
            data_im_out => mul_im_out(133)
        );

 
    UMUL_134 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(134),
            data_im_in => first_stage_im_out(134),
            re_multiplicator => re_multiplicator(134), ---  0.956970214844
            im_multiplicator => im_multiplicator(134), --- j-0.290283203125
            data_re_out => mul_re_out(134),
            data_im_out => mul_im_out(134)
        );

 
    UMUL_135 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(135),
            data_im_in => first_stage_im_out(135),
            re_multiplicator => re_multiplicator(135), ---  0.941528320312
            im_multiplicator => im_multiplicator(135), --- j-0.3369140625
            data_re_out => mul_re_out(135),
            data_im_out => mul_im_out(135)
        );

 
    UMUL_136 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(136),
            data_im_in => first_stage_im_out(136),
            re_multiplicator => re_multiplicator(136), ---  0.923889160156
            im_multiplicator => im_multiplicator(136), --- j-0.382690429688
            data_re_out => mul_re_out(136),
            data_im_out => mul_im_out(136)
        );

 
    UMUL_137 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(137),
            data_im_in => first_stage_im_out(137),
            re_multiplicator => re_multiplicator(137), ---  0.903991699219
            im_multiplicator => im_multiplicator(137), --- j-0.427551269531
            data_re_out => mul_re_out(137),
            data_im_out => mul_im_out(137)
        );

 
    UMUL_138 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(138),
            data_im_in => first_stage_im_out(138),
            re_multiplicator => re_multiplicator(138), ---  0.881896972656
            im_multiplicator => im_multiplicator(138), --- j-0.471374511719
            data_re_out => mul_re_out(138),
            data_im_out => mul_im_out(138)
        );

 
    UMUL_139 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(139),
            data_im_in => first_stage_im_out(139),
            re_multiplicator => re_multiplicator(139), ---  0.857727050781
            im_multiplicator => im_multiplicator(139), --- j-0.514099121094
            data_re_out => mul_re_out(139),
            data_im_out => mul_im_out(139)
        );

 
    UMUL_140 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(140),
            data_im_in => first_stage_im_out(140),
            re_multiplicator => re_multiplicator(140), ---  0.831481933594
            im_multiplicator => im_multiplicator(140), --- j-0.555541992188
            data_re_out => mul_re_out(140),
            data_im_out => mul_im_out(140)
        );

 
    UMUL_141 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(141),
            data_im_in => first_stage_im_out(141),
            re_multiplicator => re_multiplicator(141), ---  0.80322265625
            im_multiplicator => im_multiplicator(141), --- j-0.595703125
            data_re_out => mul_re_out(141),
            data_im_out => mul_im_out(141)
        );

 
    UMUL_142 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(142),
            data_im_in => first_stage_im_out(142),
            re_multiplicator => re_multiplicator(142), ---  0.773010253906
            im_multiplicator => im_multiplicator(142), --- j-0.634399414062
            data_re_out => mul_re_out(142),
            data_im_out => mul_im_out(142)
        );

 
    UMUL_143 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(143),
            data_im_in => first_stage_im_out(143),
            re_multiplicator => re_multiplicator(143), ---  0.740966796875
            im_multiplicator => im_multiplicator(143), --- j-0.671569824219
            data_re_out => mul_re_out(143),
            data_im_out => mul_im_out(143)
        );

 
    UMUL_144 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(144),
            data_im_in => first_stage_im_out(144),
            re_multiplicator => re_multiplicator(144), ---  0.707092285156
            im_multiplicator => im_multiplicator(144), --- j-0.707092285156
            data_re_out => mul_re_out(144),
            data_im_out => mul_im_out(144)
        );

 
    UMUL_145 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(145),
            data_im_in => first_stage_im_out(145),
            re_multiplicator => re_multiplicator(145), ---  0.671569824219
            im_multiplicator => im_multiplicator(145), --- j-0.740966796875
            data_re_out => mul_re_out(145),
            data_im_out => mul_im_out(145)
        );

 
    UMUL_146 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(146),
            data_im_in => first_stage_im_out(146),
            re_multiplicator => re_multiplicator(146), ---  0.634399414062
            im_multiplicator => im_multiplicator(146), --- j-0.773010253906
            data_re_out => mul_re_out(146),
            data_im_out => mul_im_out(146)
        );

 
    UMUL_147 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(147),
            data_im_in => first_stage_im_out(147),
            re_multiplicator => re_multiplicator(147), ---  0.595703125
            im_multiplicator => im_multiplicator(147), --- j-0.80322265625
            data_re_out => mul_re_out(147),
            data_im_out => mul_im_out(147)
        );

 
    UMUL_148 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(148),
            data_im_in => first_stage_im_out(148),
            re_multiplicator => re_multiplicator(148), ---  0.555541992188
            im_multiplicator => im_multiplicator(148), --- j-0.831481933594
            data_re_out => mul_re_out(148),
            data_im_out => mul_im_out(148)
        );

 
    UMUL_149 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(149),
            data_im_in => first_stage_im_out(149),
            re_multiplicator => re_multiplicator(149), ---  0.514099121094
            im_multiplicator => im_multiplicator(149), --- j-0.857727050781
            data_re_out => mul_re_out(149),
            data_im_out => mul_im_out(149)
        );

 
    UMUL_150 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(150),
            data_im_in => first_stage_im_out(150),
            re_multiplicator => re_multiplicator(150), ---  0.471374511719
            im_multiplicator => im_multiplicator(150), --- j-0.881896972656
            data_re_out => mul_re_out(150),
            data_im_out => mul_im_out(150)
        );

 
    UMUL_151 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(151),
            data_im_in => first_stage_im_out(151),
            re_multiplicator => re_multiplicator(151), ---  0.427551269531
            im_multiplicator => im_multiplicator(151), --- j-0.903991699219
            data_re_out => mul_re_out(151),
            data_im_out => mul_im_out(151)
        );

 
    UMUL_152 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(152),
            data_im_in => first_stage_im_out(152),
            re_multiplicator => re_multiplicator(152), ---  0.382690429688
            im_multiplicator => im_multiplicator(152), --- j-0.923889160156
            data_re_out => mul_re_out(152),
            data_im_out => mul_im_out(152)
        );

 
    UMUL_153 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(153),
            data_im_in => first_stage_im_out(153),
            re_multiplicator => re_multiplicator(153), ---  0.3369140625
            im_multiplicator => im_multiplicator(153), --- j-0.941528320312
            data_re_out => mul_re_out(153),
            data_im_out => mul_im_out(153)
        );

 
    UMUL_154 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(154),
            data_im_in => first_stage_im_out(154),
            re_multiplicator => re_multiplicator(154), ---  0.290283203125
            im_multiplicator => im_multiplicator(154), --- j-0.956970214844
            data_re_out => mul_re_out(154),
            data_im_out => mul_im_out(154)
        );

 
    UMUL_155 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(155),
            data_im_in => first_stage_im_out(155),
            re_multiplicator => re_multiplicator(155), ---  0.242980957031
            im_multiplicator => im_multiplicator(155), --- j-0.970031738281
            data_re_out => mul_re_out(155),
            data_im_out => mul_im_out(155)
        );

 
    UMUL_156 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(156),
            data_im_in => first_stage_im_out(156),
            re_multiplicator => re_multiplicator(156), ---  0.195068359375
            im_multiplicator => im_multiplicator(156), --- j-0.980773925781
            data_re_out => mul_re_out(156),
            data_im_out => mul_im_out(156)
        );

 
    UMUL_157 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(157),
            data_im_in => first_stage_im_out(157),
            re_multiplicator => re_multiplicator(157), ---  0.146728515625
            im_multiplicator => im_multiplicator(157), --- j-0.989196777344
            data_re_out => mul_re_out(157),
            data_im_out => mul_im_out(157)
        );

 
    UMUL_158 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(158),
            data_im_in => first_stage_im_out(158),
            re_multiplicator => re_multiplicator(158), ---  0.0980224609375
            im_multiplicator => im_multiplicator(158), --- j-0.995178222656
            data_re_out => mul_re_out(158),
            data_im_out => mul_im_out(158)
        );

 
    UMUL_159 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(159),
            data_im_in => first_stage_im_out(159),
            re_multiplicator => re_multiplicator(159), ---  0.049072265625
            im_multiplicator => im_multiplicator(159), --- j-0.998779296875
            data_re_out => mul_re_out(159),
            data_im_out => mul_im_out(159)
        );

 
    UMUL_160 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(160),
            data_im_in => first_stage_im_out(160),
            data_re_out => mul_re_out(160),
            data_im_out => mul_im_out(160)
        );

 
    UMUL_161 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(161),
            data_im_in => first_stage_im_out(161),
            re_multiplicator => re_multiplicator(161), ---  0.998107910156
            im_multiplicator => im_multiplicator(161), --- j-0.0613403320312
            data_re_out => mul_re_out(161),
            data_im_out => mul_im_out(161)
        );

 
    UMUL_162 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(162),
            data_im_in => first_stage_im_out(162),
            re_multiplicator => re_multiplicator(162), ---  0.992492675781
            im_multiplicator => im_multiplicator(162), --- j-0.122436523438
            data_re_out => mul_re_out(162),
            data_im_out => mul_im_out(162)
        );

 
    UMUL_163 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(163),
            data_im_in => first_stage_im_out(163),
            re_multiplicator => re_multiplicator(163), ---  0.983093261719
            im_multiplicator => im_multiplicator(163), --- j-0.183044433594
            data_re_out => mul_re_out(163),
            data_im_out => mul_im_out(163)
        );

 
    UMUL_164 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(164),
            data_im_in => first_stage_im_out(164),
            re_multiplicator => re_multiplicator(164), ---  0.970031738281
            im_multiplicator => im_multiplicator(164), --- j-0.242980957031
            data_re_out => mul_re_out(164),
            data_im_out => mul_im_out(164)
        );

 
    UMUL_165 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(165),
            data_im_in => first_stage_im_out(165),
            re_multiplicator => re_multiplicator(165), ---  0.953308105469
            im_multiplicator => im_multiplicator(165), --- j-0.302001953125
            data_re_out => mul_re_out(165),
            data_im_out => mul_im_out(165)
        );

 
    UMUL_166 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(166),
            data_im_in => first_stage_im_out(166),
            re_multiplicator => re_multiplicator(166), ---  0.932983398438
            im_multiplicator => im_multiplicator(166), --- j-0.359924316406
            data_re_out => mul_re_out(166),
            data_im_out => mul_im_out(166)
        );

 
    UMUL_167 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(167),
            data_im_in => first_stage_im_out(167),
            re_multiplicator => re_multiplicator(167), ---  0.9091796875
            im_multiplicator => im_multiplicator(167), --- j-0.416442871094
            data_re_out => mul_re_out(167),
            data_im_out => mul_im_out(167)
        );

 
    UMUL_168 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(168),
            data_im_in => first_stage_im_out(168),
            re_multiplicator => re_multiplicator(168), ---  0.881896972656
            im_multiplicator => im_multiplicator(168), --- j-0.471374511719
            data_re_out => mul_re_out(168),
            data_im_out => mul_im_out(168)
        );

 
    UMUL_169 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(169),
            data_im_in => first_stage_im_out(169),
            re_multiplicator => re_multiplicator(169), ---  0.851379394531
            im_multiplicator => im_multiplicator(169), --- j-0.524597167969
            data_re_out => mul_re_out(169),
            data_im_out => mul_im_out(169)
        );

 
    UMUL_170 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(170),
            data_im_in => first_stage_im_out(170),
            re_multiplicator => re_multiplicator(170), ---  0.817565917969
            im_multiplicator => im_multiplicator(170), --- j-0.575805664062
            data_re_out => mul_re_out(170),
            data_im_out => mul_im_out(170)
        );

 
    UMUL_171 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(171),
            data_im_in => first_stage_im_out(171),
            re_multiplicator => re_multiplicator(171), ---  0.78076171875
            im_multiplicator => im_multiplicator(171), --- j-0.624877929688
            data_re_out => mul_re_out(171),
            data_im_out => mul_im_out(171)
        );

 
    UMUL_172 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(172),
            data_im_in => first_stage_im_out(172),
            re_multiplicator => re_multiplicator(172), ---  0.740966796875
            im_multiplicator => im_multiplicator(172), --- j-0.671569824219
            data_re_out => mul_re_out(172),
            data_im_out => mul_im_out(172)
        );

 
    UMUL_173 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(173),
            data_im_in => first_stage_im_out(173),
            re_multiplicator => re_multiplicator(173), ---  0.698364257812
            im_multiplicator => im_multiplicator(173), --- j-0.715759277344
            data_re_out => mul_re_out(173),
            data_im_out => mul_im_out(173)
        );

 
    UMUL_174 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(174),
            data_im_in => first_stage_im_out(174),
            re_multiplicator => re_multiplicator(174), ---  0.653198242188
            im_multiplicator => im_multiplicator(174), --- j-0.757202148438
            data_re_out => mul_re_out(174),
            data_im_out => mul_im_out(174)
        );

 
    UMUL_175 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(175),
            data_im_in => first_stage_im_out(175),
            re_multiplicator => re_multiplicator(175), ---  0.605529785156
            im_multiplicator => im_multiplicator(175), --- j-0.795837402344
            data_re_out => mul_re_out(175),
            data_im_out => mul_im_out(175)
        );

 
    UMUL_176 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(176),
            data_im_in => first_stage_im_out(176),
            re_multiplicator => re_multiplicator(176), ---  0.555541992188
            im_multiplicator => im_multiplicator(176), --- j-0.831481933594
            data_re_out => mul_re_out(176),
            data_im_out => mul_im_out(176)
        );

 
    UMUL_177 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(177),
            data_im_in => first_stage_im_out(177),
            re_multiplicator => re_multiplicator(177), ---  0.503540039062
            im_multiplicator => im_multiplicator(177), --- j-0.863952636719
            data_re_out => mul_re_out(177),
            data_im_out => mul_im_out(177)
        );

 
    UMUL_178 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(178),
            data_im_in => first_stage_im_out(178),
            re_multiplicator => re_multiplicator(178), ---  0.449584960938
            im_multiplicator => im_multiplicator(178), --- j-0.893249511719
            data_re_out => mul_re_out(178),
            data_im_out => mul_im_out(178)
        );

 
    UMUL_179 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(179),
            data_im_in => first_stage_im_out(179),
            re_multiplicator => re_multiplicator(179), ---  0.393981933594
            im_multiplicator => im_multiplicator(179), --- j-0.919128417969
            data_re_out => mul_re_out(179),
            data_im_out => mul_im_out(179)
        );

 
    UMUL_180 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(180),
            data_im_in => first_stage_im_out(180),
            re_multiplicator => re_multiplicator(180), ---  0.3369140625
            im_multiplicator => im_multiplicator(180), --- j-0.941528320312
            data_re_out => mul_re_out(180),
            data_im_out => mul_im_out(180)
        );

 
    UMUL_181 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(181),
            data_im_in => first_stage_im_out(181),
            re_multiplicator => re_multiplicator(181), ---  0.278503417969
            im_multiplicator => im_multiplicator(181), --- j-0.96044921875
            data_re_out => mul_re_out(181),
            data_im_out => mul_im_out(181)
        );

 
    UMUL_182 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(182),
            data_im_in => first_stage_im_out(182),
            re_multiplicator => re_multiplicator(182), ---  0.219116210938
            im_multiplicator => im_multiplicator(182), --- j-0.975708007812
            data_re_out => mul_re_out(182),
            data_im_out => mul_im_out(182)
        );

 
    UMUL_183 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(183),
            data_im_in => first_stage_im_out(183),
            re_multiplicator => re_multiplicator(183), ---  0.158874511719
            im_multiplicator => im_multiplicator(183), --- j-0.9873046875
            data_re_out => mul_re_out(183),
            data_im_out => mul_im_out(183)
        );

 
    UMUL_184 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(184),
            data_im_in => first_stage_im_out(184),
            re_multiplicator => re_multiplicator(184), ---  0.0980224609375
            im_multiplicator => im_multiplicator(184), --- j-0.995178222656
            data_re_out => mul_re_out(184),
            data_im_out => mul_im_out(184)
        );

 
    UMUL_185 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(185),
            data_im_in => first_stage_im_out(185),
            re_multiplicator => re_multiplicator(185), ---  0.0368041992188
            im_multiplicator => im_multiplicator(185), --- j-0.999328613281
            data_re_out => mul_re_out(185),
            data_im_out => mul_im_out(185)
        );

 
    UMUL_186 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(186),
            data_im_in => first_stage_im_out(186),
            re_multiplicator => re_multiplicator(186), ---  -0.0245361328125
            im_multiplicator => im_multiplicator(186), --- j-0.999694824219
            data_re_out => mul_re_out(186),
            data_im_out => mul_im_out(186)
        );

 
    UMUL_187 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(187),
            data_im_in => first_stage_im_out(187),
            re_multiplicator => re_multiplicator(187), ---  -0.0858154296875
            im_multiplicator => im_multiplicator(187), --- j-0.996337890625
            data_re_out => mul_re_out(187),
            data_im_out => mul_im_out(187)
        );

 
    UMUL_188 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(188),
            data_im_in => first_stage_im_out(188),
            re_multiplicator => re_multiplicator(188), ---  -0.146728515625
            im_multiplicator => im_multiplicator(188), --- j-0.989196777344
            data_re_out => mul_re_out(188),
            data_im_out => mul_im_out(188)
        );

 
    UMUL_189 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(189),
            data_im_in => first_stage_im_out(189),
            re_multiplicator => re_multiplicator(189), ---  -0.207092285156
            im_multiplicator => im_multiplicator(189), --- j-0.978332519531
            data_re_out => mul_re_out(189),
            data_im_out => mul_im_out(189)
        );

 
    UMUL_190 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(190),
            data_im_in => first_stage_im_out(190),
            re_multiplicator => re_multiplicator(190), ---  -0.266723632812
            im_multiplicator => im_multiplicator(190), --- j-0.963806152344
            data_re_out => mul_re_out(190),
            data_im_out => mul_im_out(190)
        );

 
    UMUL_191 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(191),
            data_im_in => first_stage_im_out(191),
            re_multiplicator => re_multiplicator(191), ---  -0.325317382812
            im_multiplicator => im_multiplicator(191), --- j-0.945617675781
            data_re_out => mul_re_out(191),
            data_im_out => mul_im_out(191)
        );

 
    UMUL_192 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(192),
            data_im_in => first_stage_im_out(192),
            data_re_out => mul_re_out(192),
            data_im_out => mul_im_out(192)
        );

 
    UMUL_193 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(193),
            data_im_in => first_stage_im_out(193),
            re_multiplicator => re_multiplicator(193), ---  0.997314453125
            im_multiplicator => im_multiplicator(193), --- j-0.0735473632812
            data_re_out => mul_re_out(193),
            data_im_out => mul_im_out(193)
        );

 
    UMUL_194 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(194),
            data_im_in => first_stage_im_out(194),
            re_multiplicator => re_multiplicator(194), ---  0.989196777344
            im_multiplicator => im_multiplicator(194), --- j-0.146728515625
            data_re_out => mul_re_out(194),
            data_im_out => mul_im_out(194)
        );

 
    UMUL_195 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(195),
            data_im_in => first_stage_im_out(195),
            re_multiplicator => re_multiplicator(195), ---  0.975708007812
            im_multiplicator => im_multiplicator(195), --- j-0.219116210938
            data_re_out => mul_re_out(195),
            data_im_out => mul_im_out(195)
        );

 
    UMUL_196 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(196),
            data_im_in => first_stage_im_out(196),
            re_multiplicator => re_multiplicator(196), ---  0.956970214844
            im_multiplicator => im_multiplicator(196), --- j-0.290283203125
            data_re_out => mul_re_out(196),
            data_im_out => mul_im_out(196)
        );

 
    UMUL_197 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(197),
            data_im_in => first_stage_im_out(197),
            re_multiplicator => re_multiplicator(197), ---  0.932983398438
            im_multiplicator => im_multiplicator(197), --- j-0.359924316406
            data_re_out => mul_re_out(197),
            data_im_out => mul_im_out(197)
        );

 
    UMUL_198 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(198),
            data_im_in => first_stage_im_out(198),
            re_multiplicator => re_multiplicator(198), ---  0.903991699219
            im_multiplicator => im_multiplicator(198), --- j-0.427551269531
            data_re_out => mul_re_out(198),
            data_im_out => mul_im_out(198)
        );

 
    UMUL_199 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(199),
            data_im_in => first_stage_im_out(199),
            re_multiplicator => re_multiplicator(199), ---  0.8701171875
            im_multiplicator => im_multiplicator(199), --- j-0.492919921875
            data_re_out => mul_re_out(199),
            data_im_out => mul_im_out(199)
        );

 
    UMUL_200 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(200),
            data_im_in => first_stage_im_out(200),
            re_multiplicator => re_multiplicator(200), ---  0.831481933594
            im_multiplicator => im_multiplicator(200), --- j-0.555541992188
            data_re_out => mul_re_out(200),
            data_im_out => mul_im_out(200)
        );

 
    UMUL_201 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(201),
            data_im_in => first_stage_im_out(201),
            re_multiplicator => re_multiplicator(201), ---  0.788330078125
            im_multiplicator => im_multiplicator(201), --- j-0.615234375
            data_re_out => mul_re_out(201),
            data_im_out => mul_im_out(201)
        );

 
    UMUL_202 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(202),
            data_im_in => first_stage_im_out(202),
            re_multiplicator => re_multiplicator(202), ---  0.740966796875
            im_multiplicator => im_multiplicator(202), --- j-0.671569824219
            data_re_out => mul_re_out(202),
            data_im_out => mul_im_out(202)
        );

 
    UMUL_203 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(203),
            data_im_in => first_stage_im_out(203),
            re_multiplicator => re_multiplicator(203), ---  0.689514160156
            im_multiplicator => im_multiplicator(203), --- j-0.724243164062
            data_re_out => mul_re_out(203),
            data_im_out => mul_im_out(203)
        );

 
    UMUL_204 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(204),
            data_im_in => first_stage_im_out(204),
            re_multiplicator => re_multiplicator(204), ---  0.634399414062
            im_multiplicator => im_multiplicator(204), --- j-0.773010253906
            data_re_out => mul_re_out(204),
            data_im_out => mul_im_out(204)
        );

 
    UMUL_205 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(205),
            data_im_in => first_stage_im_out(205),
            re_multiplicator => re_multiplicator(205), ---  0.575805664062
            im_multiplicator => im_multiplicator(205), --- j-0.817565917969
            data_re_out => mul_re_out(205),
            data_im_out => mul_im_out(205)
        );

 
    UMUL_206 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(206),
            data_im_in => first_stage_im_out(206),
            re_multiplicator => re_multiplicator(206), ---  0.514099121094
            im_multiplicator => im_multiplicator(206), --- j-0.857727050781
            data_re_out => mul_re_out(206),
            data_im_out => mul_im_out(206)
        );

 
    UMUL_207 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(207),
            data_im_in => first_stage_im_out(207),
            re_multiplicator => re_multiplicator(207), ---  0.449584960938
            im_multiplicator => im_multiplicator(207), --- j-0.893249511719
            data_re_out => mul_re_out(207),
            data_im_out => mul_im_out(207)
        );

 
    UMUL_208 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(208),
            data_im_in => first_stage_im_out(208),
            re_multiplicator => re_multiplicator(208), ---  0.382690429688
            im_multiplicator => im_multiplicator(208), --- j-0.923889160156
            data_re_out => mul_re_out(208),
            data_im_out => mul_im_out(208)
        );

 
    UMUL_209 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(209),
            data_im_in => first_stage_im_out(209),
            re_multiplicator => re_multiplicator(209), ---  0.313659667969
            im_multiplicator => im_multiplicator(209), --- j-0.949523925781
            data_re_out => mul_re_out(209),
            data_im_out => mul_im_out(209)
        );

 
    UMUL_210 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(210),
            data_im_in => first_stage_im_out(210),
            re_multiplicator => re_multiplicator(210), ---  0.242980957031
            im_multiplicator => im_multiplicator(210), --- j-0.970031738281
            data_re_out => mul_re_out(210),
            data_im_out => mul_im_out(210)
        );

 
    UMUL_211 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(211),
            data_im_in => first_stage_im_out(211),
            re_multiplicator => re_multiplicator(211), ---  0.170959472656
            im_multiplicator => im_multiplicator(211), --- j-0.985290527344
            data_re_out => mul_re_out(211),
            data_im_out => mul_im_out(211)
        );

 
    UMUL_212 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(212),
            data_im_in => first_stage_im_out(212),
            re_multiplicator => re_multiplicator(212), ---  0.0980224609375
            im_multiplicator => im_multiplicator(212), --- j-0.995178222656
            data_re_out => mul_re_out(212),
            data_im_out => mul_im_out(212)
        );

 
    UMUL_213 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(213),
            data_im_in => first_stage_im_out(213),
            re_multiplicator => re_multiplicator(213), ---  0.0245361328125
            im_multiplicator => im_multiplicator(213), --- j-0.999694824219
            data_re_out => mul_re_out(213),
            data_im_out => mul_im_out(213)
        );

 
    UMUL_214 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(214),
            data_im_in => first_stage_im_out(214),
            re_multiplicator => re_multiplicator(214), ---  -0.049072265625
            im_multiplicator => im_multiplicator(214), --- j-0.998779296875
            data_re_out => mul_re_out(214),
            data_im_out => mul_im_out(214)
        );

 
    UMUL_215 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(215),
            data_im_in => first_stage_im_out(215),
            re_multiplicator => re_multiplicator(215), ---  -0.122436523438
            im_multiplicator => im_multiplicator(215), --- j-0.992492675781
            data_re_out => mul_re_out(215),
            data_im_out => mul_im_out(215)
        );

 
    UMUL_216 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(216),
            data_im_in => first_stage_im_out(216),
            re_multiplicator => re_multiplicator(216), ---  -0.195068359375
            im_multiplicator => im_multiplicator(216), --- j-0.980773925781
            data_re_out => mul_re_out(216),
            data_im_out => mul_im_out(216)
        );

 
    UMUL_217 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(217),
            data_im_in => first_stage_im_out(217),
            re_multiplicator => re_multiplicator(217), ---  -0.266723632812
            im_multiplicator => im_multiplicator(217), --- j-0.963806152344
            data_re_out => mul_re_out(217),
            data_im_out => mul_im_out(217)
        );

 
    UMUL_218 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(218),
            data_im_in => first_stage_im_out(218),
            re_multiplicator => re_multiplicator(218), ---  -0.3369140625
            im_multiplicator => im_multiplicator(218), --- j-0.941528320312
            data_re_out => mul_re_out(218),
            data_im_out => mul_im_out(218)
        );

 
    UMUL_219 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(219),
            data_im_in => first_stage_im_out(219),
            re_multiplicator => re_multiplicator(219), ---  -0.405212402344
            im_multiplicator => im_multiplicator(219), --- j-0.914184570312
            data_re_out => mul_re_out(219),
            data_im_out => mul_im_out(219)
        );

 
    UMUL_220 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(220),
            data_im_in => first_stage_im_out(220),
            re_multiplicator => re_multiplicator(220), ---  -0.471374511719
            im_multiplicator => im_multiplicator(220), --- j-0.881896972656
            data_re_out => mul_re_out(220),
            data_im_out => mul_im_out(220)
        );

 
    UMUL_221 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(221),
            data_im_in => first_stage_im_out(221),
            re_multiplicator => re_multiplicator(221), ---  -0.534973144531
            im_multiplicator => im_multiplicator(221), --- j-0.844848632812
            data_re_out => mul_re_out(221),
            data_im_out => mul_im_out(221)
        );

 
    UMUL_222 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(222),
            data_im_in => first_stage_im_out(222),
            re_multiplicator => re_multiplicator(222), ---  -0.595703125
            im_multiplicator => im_multiplicator(222), --- j-0.80322265625
            data_re_out => mul_re_out(222),
            data_im_out => mul_im_out(222)
        );

 
    UMUL_223 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(223),
            data_im_in => first_stage_im_out(223),
            re_multiplicator => re_multiplicator(223), ---  -0.653198242188
            im_multiplicator => im_multiplicator(223), --- j-0.757202148438
            data_re_out => mul_re_out(223),
            data_im_out => mul_im_out(223)
        );

 
    UMUL_224 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(224),
            data_im_in => first_stage_im_out(224),
            data_re_out => mul_re_out(224),
            data_im_out => mul_im_out(224)
        );

 
    UMUL_225 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(225),
            data_im_in => first_stage_im_out(225),
            re_multiplicator => re_multiplicator(225), ---  0.996337890625
            im_multiplicator => im_multiplicator(225), --- j-0.0858154296875
            data_re_out => mul_re_out(225),
            data_im_out => mul_im_out(225)
        );

 
    UMUL_226 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(226),
            data_im_in => first_stage_im_out(226),
            re_multiplicator => re_multiplicator(226), ---  0.985290527344
            im_multiplicator => im_multiplicator(226), --- j-0.170959472656
            data_re_out => mul_re_out(226),
            data_im_out => mul_im_out(226)
        );

 
    UMUL_227 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(227),
            data_im_in => first_stage_im_out(227),
            re_multiplicator => re_multiplicator(227), ---  0.966979980469
            im_multiplicator => im_multiplicator(227), --- j-0.2548828125
            data_re_out => mul_re_out(227),
            data_im_out => mul_im_out(227)
        );

 
    UMUL_228 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(228),
            data_im_in => first_stage_im_out(228),
            re_multiplicator => re_multiplicator(228), ---  0.941528320312
            im_multiplicator => im_multiplicator(228), --- j-0.3369140625
            data_re_out => mul_re_out(228),
            data_im_out => mul_im_out(228)
        );

 
    UMUL_229 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(229),
            data_im_in => first_stage_im_out(229),
            re_multiplicator => re_multiplicator(229), ---  0.9091796875
            im_multiplicator => im_multiplicator(229), --- j-0.416442871094
            data_re_out => mul_re_out(229),
            data_im_out => mul_im_out(229)
        );

 
    UMUL_230 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(230),
            data_im_in => first_stage_im_out(230),
            re_multiplicator => re_multiplicator(230), ---  0.8701171875
            im_multiplicator => im_multiplicator(230), --- j-0.492919921875
            data_re_out => mul_re_out(230),
            data_im_out => mul_im_out(230)
        );

 
    UMUL_231 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(231),
            data_im_in => first_stage_im_out(231),
            re_multiplicator => re_multiplicator(231), ---  0.824584960938
            im_multiplicator => im_multiplicator(231), --- j-0.565734863281
            data_re_out => mul_re_out(231),
            data_im_out => mul_im_out(231)
        );

 
    UMUL_232 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(232),
            data_im_in => first_stage_im_out(232),
            re_multiplicator => re_multiplicator(232), ---  0.773010253906
            im_multiplicator => im_multiplicator(232), --- j-0.634399414062
            data_re_out => mul_re_out(232),
            data_im_out => mul_im_out(232)
        );

 
    UMUL_233 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(233),
            data_im_in => first_stage_im_out(233),
            re_multiplicator => re_multiplicator(233), ---  0.715759277344
            im_multiplicator => im_multiplicator(233), --- j-0.698364257812
            data_re_out => mul_re_out(233),
            data_im_out => mul_im_out(233)
        );

 
    UMUL_234 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(234),
            data_im_in => first_stage_im_out(234),
            re_multiplicator => re_multiplicator(234), ---  0.653198242188
            im_multiplicator => im_multiplicator(234), --- j-0.757202148438
            data_re_out => mul_re_out(234),
            data_im_out => mul_im_out(234)
        );

 
    UMUL_235 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(235),
            data_im_in => first_stage_im_out(235),
            re_multiplicator => re_multiplicator(235), ---  0.585815429688
            im_multiplicator => im_multiplicator(235), --- j-0.810485839844
            data_re_out => mul_re_out(235),
            data_im_out => mul_im_out(235)
        );

 
    UMUL_236 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(236),
            data_im_in => first_stage_im_out(236),
            re_multiplicator => re_multiplicator(236), ---  0.514099121094
            im_multiplicator => im_multiplicator(236), --- j-0.857727050781
            data_re_out => mul_re_out(236),
            data_im_out => mul_im_out(236)
        );

 
    UMUL_237 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(237),
            data_im_in => first_stage_im_out(237),
            re_multiplicator => re_multiplicator(237), ---  0.438598632812
            im_multiplicator => im_multiplicator(237), --- j-0.898681640625
            data_re_out => mul_re_out(237),
            data_im_out => mul_im_out(237)
        );

 
    UMUL_238 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(238),
            data_im_in => first_stage_im_out(238),
            re_multiplicator => re_multiplicator(238), ---  0.359924316406
            im_multiplicator => im_multiplicator(238), --- j-0.932983398438
            data_re_out => mul_re_out(238),
            data_im_out => mul_im_out(238)
        );

 
    UMUL_239 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(239),
            data_im_in => first_stage_im_out(239),
            re_multiplicator => re_multiplicator(239), ---  0.278503417969
            im_multiplicator => im_multiplicator(239), --- j-0.96044921875
            data_re_out => mul_re_out(239),
            data_im_out => mul_im_out(239)
        );

 
    UMUL_240 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(240),
            data_im_in => first_stage_im_out(240),
            re_multiplicator => re_multiplicator(240), ---  0.195068359375
            im_multiplicator => im_multiplicator(240), --- j-0.980773925781
            data_re_out => mul_re_out(240),
            data_im_out => mul_im_out(240)
        );

 
    UMUL_241 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(241),
            data_im_in => first_stage_im_out(241),
            re_multiplicator => re_multiplicator(241), ---  0.110229492188
            im_multiplicator => im_multiplicator(241), --- j-0.993896484375
            data_re_out => mul_re_out(241),
            data_im_out => mul_im_out(241)
        );

 
    UMUL_242 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(242),
            data_im_in => first_stage_im_out(242),
            re_multiplicator => re_multiplicator(242), ---  0.0245361328125
            im_multiplicator => im_multiplicator(242), --- j-0.999694824219
            data_re_out => mul_re_out(242),
            data_im_out => mul_im_out(242)
        );

 
    UMUL_243 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(243),
            data_im_in => first_stage_im_out(243),
            re_multiplicator => re_multiplicator(243), ---  -0.0613403320312
            im_multiplicator => im_multiplicator(243), --- j-0.998107910156
            data_re_out => mul_re_out(243),
            data_im_out => mul_im_out(243)
        );

 
    UMUL_244 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(244),
            data_im_in => first_stage_im_out(244),
            re_multiplicator => re_multiplicator(244), ---  -0.146728515625
            im_multiplicator => im_multiplicator(244), --- j-0.989196777344
            data_re_out => mul_re_out(244),
            data_im_out => mul_im_out(244)
        );

 
    UMUL_245 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(245),
            data_im_in => first_stage_im_out(245),
            re_multiplicator => re_multiplicator(245), ---  -0.231079101562
            im_multiplicator => im_multiplicator(245), --- j-0.972961425781
            data_re_out => mul_re_out(245),
            data_im_out => mul_im_out(245)
        );

 
    UMUL_246 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(246),
            data_im_in => first_stage_im_out(246),
            re_multiplicator => re_multiplicator(246), ---  -0.313659667969
            im_multiplicator => im_multiplicator(246), --- j-0.949523925781
            data_re_out => mul_re_out(246),
            data_im_out => mul_im_out(246)
        );

 
    UMUL_247 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(247),
            data_im_in => first_stage_im_out(247),
            re_multiplicator => re_multiplicator(247), ---  -0.393981933594
            im_multiplicator => im_multiplicator(247), --- j-0.919128417969
            data_re_out => mul_re_out(247),
            data_im_out => mul_im_out(247)
        );

 
    UMUL_248 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(248),
            data_im_in => first_stage_im_out(248),
            re_multiplicator => re_multiplicator(248), ---  -0.471374511719
            im_multiplicator => im_multiplicator(248), --- j-0.881896972656
            data_re_out => mul_re_out(248),
            data_im_out => mul_im_out(248)
        );

 
    UMUL_249 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(249),
            data_im_in => first_stage_im_out(249),
            re_multiplicator => re_multiplicator(249), ---  -0.545349121094
            im_multiplicator => im_multiplicator(249), --- j-0.838195800781
            data_re_out => mul_re_out(249),
            data_im_out => mul_im_out(249)
        );

 
    UMUL_250 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(250),
            data_im_in => first_stage_im_out(250),
            re_multiplicator => re_multiplicator(250), ---  -0.615234375
            im_multiplicator => im_multiplicator(250), --- j-0.788330078125
            data_re_out => mul_re_out(250),
            data_im_out => mul_im_out(250)
        );

 
    UMUL_251 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(251),
            data_im_in => first_stage_im_out(251),
            re_multiplicator => re_multiplicator(251), ---  -0.680603027344
            im_multiplicator => im_multiplicator(251), --- j-0.732666015625
            data_re_out => mul_re_out(251),
            data_im_out => mul_im_out(251)
        );

 
    UMUL_252 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(252),
            data_im_in => first_stage_im_out(252),
            re_multiplicator => re_multiplicator(252), ---  -0.740966796875
            im_multiplicator => im_multiplicator(252), --- j-0.671569824219
            data_re_out => mul_re_out(252),
            data_im_out => mul_im_out(252)
        );

 
    UMUL_253 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(253),
            data_im_in => first_stage_im_out(253),
            re_multiplicator => re_multiplicator(253), ---  -0.795837402344
            im_multiplicator => im_multiplicator(253), --- j-0.605529785156
            data_re_out => mul_re_out(253),
            data_im_out => mul_im_out(253)
        );

 
    UMUL_254 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(254),
            data_im_in => first_stage_im_out(254),
            re_multiplicator => re_multiplicator(254), ---  -0.844848632812
            im_multiplicator => im_multiplicator(254), --- j-0.534973144531
            data_re_out => mul_re_out(254),
            data_im_out => mul_im_out(254)
        );

 
    UMUL_255 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(255),
            data_im_in => first_stage_im_out(255),
            re_multiplicator => re_multiplicator(255), ---  -0.887634277344
            im_multiplicator => im_multiplicator(255), --- j-0.460510253906
            data_re_out => mul_re_out(255),
            data_im_out => mul_im_out(255)
        );

 
    UMUL_256 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(256),
            data_im_in => first_stage_im_out(256),
            data_re_out => mul_re_out(256),
            data_im_out => mul_im_out(256)
        );

 
    UMUL_257 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(257),
            data_im_in => first_stage_im_out(257),
            re_multiplicator => re_multiplicator(257), ---  0.995178222656
            im_multiplicator => im_multiplicator(257), --- j-0.0980224609375
            data_re_out => mul_re_out(257),
            data_im_out => mul_im_out(257)
        );

 
    UMUL_258 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(258),
            data_im_in => first_stage_im_out(258),
            re_multiplicator => re_multiplicator(258), ---  0.980773925781
            im_multiplicator => im_multiplicator(258), --- j-0.195068359375
            data_re_out => mul_re_out(258),
            data_im_out => mul_im_out(258)
        );

 
    UMUL_259 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(259),
            data_im_in => first_stage_im_out(259),
            re_multiplicator => re_multiplicator(259), ---  0.956970214844
            im_multiplicator => im_multiplicator(259), --- j-0.290283203125
            data_re_out => mul_re_out(259),
            data_im_out => mul_im_out(259)
        );

 
    UMUL_260 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(260),
            data_im_in => first_stage_im_out(260),
            re_multiplicator => re_multiplicator(260), ---  0.923889160156
            im_multiplicator => im_multiplicator(260), --- j-0.382690429688
            data_re_out => mul_re_out(260),
            data_im_out => mul_im_out(260)
        );

 
    UMUL_261 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(261),
            data_im_in => first_stage_im_out(261),
            re_multiplicator => re_multiplicator(261), ---  0.881896972656
            im_multiplicator => im_multiplicator(261), --- j-0.471374511719
            data_re_out => mul_re_out(261),
            data_im_out => mul_im_out(261)
        );

 
    UMUL_262 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(262),
            data_im_in => first_stage_im_out(262),
            re_multiplicator => re_multiplicator(262), ---  0.831481933594
            im_multiplicator => im_multiplicator(262), --- j-0.555541992188
            data_re_out => mul_re_out(262),
            data_im_out => mul_im_out(262)
        );

 
    UMUL_263 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(263),
            data_im_in => first_stage_im_out(263),
            re_multiplicator => re_multiplicator(263), ---  0.773010253906
            im_multiplicator => im_multiplicator(263), --- j-0.634399414062
            data_re_out => mul_re_out(263),
            data_im_out => mul_im_out(263)
        );

 
    UMUL_264 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(264),
            data_im_in => first_stage_im_out(264),
            re_multiplicator => re_multiplicator(264), ---  0.707092285156
            im_multiplicator => im_multiplicator(264), --- j-0.707092285156
            data_re_out => mul_re_out(264),
            data_im_out => mul_im_out(264)
        );

 
    UMUL_265 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(265),
            data_im_in => first_stage_im_out(265),
            re_multiplicator => re_multiplicator(265), ---  0.634399414062
            im_multiplicator => im_multiplicator(265), --- j-0.773010253906
            data_re_out => mul_re_out(265),
            data_im_out => mul_im_out(265)
        );

 
    UMUL_266 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(266),
            data_im_in => first_stage_im_out(266),
            re_multiplicator => re_multiplicator(266), ---  0.555541992188
            im_multiplicator => im_multiplicator(266), --- j-0.831481933594
            data_re_out => mul_re_out(266),
            data_im_out => mul_im_out(266)
        );

 
    UMUL_267 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(267),
            data_im_in => first_stage_im_out(267),
            re_multiplicator => re_multiplicator(267), ---  0.471374511719
            im_multiplicator => im_multiplicator(267), --- j-0.881896972656
            data_re_out => mul_re_out(267),
            data_im_out => mul_im_out(267)
        );

 
    UMUL_268 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(268),
            data_im_in => first_stage_im_out(268),
            re_multiplicator => re_multiplicator(268), ---  0.382690429688
            im_multiplicator => im_multiplicator(268), --- j-0.923889160156
            data_re_out => mul_re_out(268),
            data_im_out => mul_im_out(268)
        );

 
    UMUL_269 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(269),
            data_im_in => first_stage_im_out(269),
            re_multiplicator => re_multiplicator(269), ---  0.290283203125
            im_multiplicator => im_multiplicator(269), --- j-0.956970214844
            data_re_out => mul_re_out(269),
            data_im_out => mul_im_out(269)
        );

 
    UMUL_270 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(270),
            data_im_in => first_stage_im_out(270),
            re_multiplicator => re_multiplicator(270), ---  0.195068359375
            im_multiplicator => im_multiplicator(270), --- j-0.980773925781
            data_re_out => mul_re_out(270),
            data_im_out => mul_im_out(270)
        );

 
    UMUL_271 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(271),
            data_im_in => first_stage_im_out(271),
            re_multiplicator => re_multiplicator(271), ---  0.0980224609375
            im_multiplicator => im_multiplicator(271), --- j-0.995178222656
            data_re_out => mul_re_out(271),
            data_im_out => mul_im_out(271)
        );

 
    UMUL_272 : multiplier_mulminusj
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(272),
            data_im_in => first_stage_im_out(272),
            data_re_out => mul_re_out(272),
            data_im_out => mul_im_out(272)
        );

 
    UMUL_273 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(273),
            data_im_in => first_stage_im_out(273),
            re_multiplicator => re_multiplicator(273), ---  -0.0980224609375
            im_multiplicator => im_multiplicator(273), --- j-0.995178222656
            data_re_out => mul_re_out(273),
            data_im_out => mul_im_out(273)
        );

 
    UMUL_274 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(274),
            data_im_in => first_stage_im_out(274),
            re_multiplicator => re_multiplicator(274), ---  -0.195068359375
            im_multiplicator => im_multiplicator(274), --- j-0.980773925781
            data_re_out => mul_re_out(274),
            data_im_out => mul_im_out(274)
        );

 
    UMUL_275 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(275),
            data_im_in => first_stage_im_out(275),
            re_multiplicator => re_multiplicator(275), ---  -0.290283203125
            im_multiplicator => im_multiplicator(275), --- j-0.956970214844
            data_re_out => mul_re_out(275),
            data_im_out => mul_im_out(275)
        );

 
    UMUL_276 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(276),
            data_im_in => first_stage_im_out(276),
            re_multiplicator => re_multiplicator(276), ---  -0.382690429688
            im_multiplicator => im_multiplicator(276), --- j-0.923889160156
            data_re_out => mul_re_out(276),
            data_im_out => mul_im_out(276)
        );

 
    UMUL_277 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(277),
            data_im_in => first_stage_im_out(277),
            re_multiplicator => re_multiplicator(277), ---  -0.471374511719
            im_multiplicator => im_multiplicator(277), --- j-0.881896972656
            data_re_out => mul_re_out(277),
            data_im_out => mul_im_out(277)
        );

 
    UMUL_278 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(278),
            data_im_in => first_stage_im_out(278),
            re_multiplicator => re_multiplicator(278), ---  -0.555541992188
            im_multiplicator => im_multiplicator(278), --- j-0.831481933594
            data_re_out => mul_re_out(278),
            data_im_out => mul_im_out(278)
        );

 
    UMUL_279 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(279),
            data_im_in => first_stage_im_out(279),
            re_multiplicator => re_multiplicator(279), ---  -0.634399414062
            im_multiplicator => im_multiplicator(279), --- j-0.773010253906
            data_re_out => mul_re_out(279),
            data_im_out => mul_im_out(279)
        );

 
    UMUL_280 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(280),
            data_im_in => first_stage_im_out(280),
            re_multiplicator => re_multiplicator(280), ---  -0.707092285156
            im_multiplicator => im_multiplicator(280), --- j-0.707092285156
            data_re_out => mul_re_out(280),
            data_im_out => mul_im_out(280)
        );

 
    UMUL_281 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(281),
            data_im_in => first_stage_im_out(281),
            re_multiplicator => re_multiplicator(281), ---  -0.773010253906
            im_multiplicator => im_multiplicator(281), --- j-0.634399414062
            data_re_out => mul_re_out(281),
            data_im_out => mul_im_out(281)
        );

 
    UMUL_282 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(282),
            data_im_in => first_stage_im_out(282),
            re_multiplicator => re_multiplicator(282), ---  -0.831481933594
            im_multiplicator => im_multiplicator(282), --- j-0.555541992188
            data_re_out => mul_re_out(282),
            data_im_out => mul_im_out(282)
        );

 
    UMUL_283 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(283),
            data_im_in => first_stage_im_out(283),
            re_multiplicator => re_multiplicator(283), ---  -0.881896972656
            im_multiplicator => im_multiplicator(283), --- j-0.471374511719
            data_re_out => mul_re_out(283),
            data_im_out => mul_im_out(283)
        );

 
    UMUL_284 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(284),
            data_im_in => first_stage_im_out(284),
            re_multiplicator => re_multiplicator(284), ---  -0.923889160156
            im_multiplicator => im_multiplicator(284), --- j-0.382690429688
            data_re_out => mul_re_out(284),
            data_im_out => mul_im_out(284)
        );

 
    UMUL_285 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(285),
            data_im_in => first_stage_im_out(285),
            re_multiplicator => re_multiplicator(285), ---  -0.956970214844
            im_multiplicator => im_multiplicator(285), --- j-0.290283203125
            data_re_out => mul_re_out(285),
            data_im_out => mul_im_out(285)
        );

 
    UMUL_286 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(286),
            data_im_in => first_stage_im_out(286),
            re_multiplicator => re_multiplicator(286), ---  -0.980773925781
            im_multiplicator => im_multiplicator(286), --- j-0.195068359375
            data_re_out => mul_re_out(286),
            data_im_out => mul_im_out(286)
        );

 
    UMUL_287 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(287),
            data_im_in => first_stage_im_out(287),
            re_multiplicator => re_multiplicator(287), ---  -0.995178222656
            im_multiplicator => im_multiplicator(287), --- j-0.0980224609375
            data_re_out => mul_re_out(287),
            data_im_out => mul_im_out(287)
        );

 
    UMUL_288 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(288),
            data_im_in => first_stage_im_out(288),
            data_re_out => mul_re_out(288),
            data_im_out => mul_im_out(288)
        );

 
    UMUL_289 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(289),
            data_im_in => first_stage_im_out(289),
            re_multiplicator => re_multiplicator(289), ---  0.993896484375
            im_multiplicator => im_multiplicator(289), --- j-0.110229492188
            data_re_out => mul_re_out(289),
            data_im_out => mul_im_out(289)
        );

 
    UMUL_290 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(290),
            data_im_in => first_stage_im_out(290),
            re_multiplicator => re_multiplicator(290), ---  0.975708007812
            im_multiplicator => im_multiplicator(290), --- j-0.219116210938
            data_re_out => mul_re_out(290),
            data_im_out => mul_im_out(290)
        );

 
    UMUL_291 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(291),
            data_im_in => first_stage_im_out(291),
            re_multiplicator => re_multiplicator(291), ---  0.945617675781
            im_multiplicator => im_multiplicator(291), --- j-0.325317382812
            data_re_out => mul_re_out(291),
            data_im_out => mul_im_out(291)
        );

 
    UMUL_292 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(292),
            data_im_in => first_stage_im_out(292),
            re_multiplicator => re_multiplicator(292), ---  0.903991699219
            im_multiplicator => im_multiplicator(292), --- j-0.427551269531
            data_re_out => mul_re_out(292),
            data_im_out => mul_im_out(292)
        );

 
    UMUL_293 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(293),
            data_im_in => first_stage_im_out(293),
            re_multiplicator => re_multiplicator(293), ---  0.851379394531
            im_multiplicator => im_multiplicator(293), --- j-0.524597167969
            data_re_out => mul_re_out(293),
            data_im_out => mul_im_out(293)
        );

 
    UMUL_294 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(294),
            data_im_in => first_stage_im_out(294),
            re_multiplicator => re_multiplicator(294), ---  0.788330078125
            im_multiplicator => im_multiplicator(294), --- j-0.615234375
            data_re_out => mul_re_out(294),
            data_im_out => mul_im_out(294)
        );

 
    UMUL_295 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(295),
            data_im_in => first_stage_im_out(295),
            re_multiplicator => re_multiplicator(295), ---  0.715759277344
            im_multiplicator => im_multiplicator(295), --- j-0.698364257812
            data_re_out => mul_re_out(295),
            data_im_out => mul_im_out(295)
        );

 
    UMUL_296 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(296),
            data_im_in => first_stage_im_out(296),
            re_multiplicator => re_multiplicator(296), ---  0.634399414062
            im_multiplicator => im_multiplicator(296), --- j-0.773010253906
            data_re_out => mul_re_out(296),
            data_im_out => mul_im_out(296)
        );

 
    UMUL_297 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(297),
            data_im_in => first_stage_im_out(297),
            re_multiplicator => re_multiplicator(297), ---  0.545349121094
            im_multiplicator => im_multiplicator(297), --- j-0.838195800781
            data_re_out => mul_re_out(297),
            data_im_out => mul_im_out(297)
        );

 
    UMUL_298 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(298),
            data_im_in => first_stage_im_out(298),
            re_multiplicator => re_multiplicator(298), ---  0.449584960938
            im_multiplicator => im_multiplicator(298), --- j-0.893249511719
            data_re_out => mul_re_out(298),
            data_im_out => mul_im_out(298)
        );

 
    UMUL_299 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(299),
            data_im_in => first_stage_im_out(299),
            re_multiplicator => re_multiplicator(299), ---  0.348388671875
            im_multiplicator => im_multiplicator(299), --- j-0.937316894531
            data_re_out => mul_re_out(299),
            data_im_out => mul_im_out(299)
        );

 
    UMUL_300 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(300),
            data_im_in => first_stage_im_out(300),
            re_multiplicator => re_multiplicator(300), ---  0.242980957031
            im_multiplicator => im_multiplicator(300), --- j-0.970031738281
            data_re_out => mul_re_out(300),
            data_im_out => mul_im_out(300)
        );

 
    UMUL_301 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(301),
            data_im_in => first_stage_im_out(301),
            re_multiplicator => re_multiplicator(301), ---  0.134582519531
            im_multiplicator => im_multiplicator(301), --- j-0.990905761719
            data_re_out => mul_re_out(301),
            data_im_out => mul_im_out(301)
        );

 
    UMUL_302 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(302),
            data_im_in => first_stage_im_out(302),
            re_multiplicator => re_multiplicator(302), ---  0.0245361328125
            im_multiplicator => im_multiplicator(302), --- j-0.999694824219
            data_re_out => mul_re_out(302),
            data_im_out => mul_im_out(302)
        );

 
    UMUL_303 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(303),
            data_im_in => first_stage_im_out(303),
            re_multiplicator => re_multiplicator(303), ---  -0.0858154296875
            im_multiplicator => im_multiplicator(303), --- j-0.996337890625
            data_re_out => mul_re_out(303),
            data_im_out => mul_im_out(303)
        );

 
    UMUL_304 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(304),
            data_im_in => first_stage_im_out(304),
            re_multiplicator => re_multiplicator(304), ---  -0.195068359375
            im_multiplicator => im_multiplicator(304), --- j-0.980773925781
            data_re_out => mul_re_out(304),
            data_im_out => mul_im_out(304)
        );

 
    UMUL_305 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(305),
            data_im_in => first_stage_im_out(305),
            re_multiplicator => re_multiplicator(305), ---  -0.302001953125
            im_multiplicator => im_multiplicator(305), --- j-0.953308105469
            data_re_out => mul_re_out(305),
            data_im_out => mul_im_out(305)
        );

 
    UMUL_306 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(306),
            data_im_in => first_stage_im_out(306),
            re_multiplicator => re_multiplicator(306), ---  -0.405212402344
            im_multiplicator => im_multiplicator(306), --- j-0.914184570312
            data_re_out => mul_re_out(306),
            data_im_out => mul_im_out(306)
        );

 
    UMUL_307 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(307),
            data_im_in => first_stage_im_out(307),
            re_multiplicator => re_multiplicator(307), ---  -0.503540039062
            im_multiplicator => im_multiplicator(307), --- j-0.863952636719
            data_re_out => mul_re_out(307),
            data_im_out => mul_im_out(307)
        );

 
    UMUL_308 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(308),
            data_im_in => first_stage_im_out(308),
            re_multiplicator => re_multiplicator(308), ---  -0.595703125
            im_multiplicator => im_multiplicator(308), --- j-0.80322265625
            data_re_out => mul_re_out(308),
            data_im_out => mul_im_out(308)
        );

 
    UMUL_309 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(309),
            data_im_in => first_stage_im_out(309),
            re_multiplicator => re_multiplicator(309), ---  -0.680603027344
            im_multiplicator => im_multiplicator(309), --- j-0.732666015625
            data_re_out => mul_re_out(309),
            data_im_out => mul_im_out(309)
        );

 
    UMUL_310 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(310),
            data_im_in => first_stage_im_out(310),
            re_multiplicator => re_multiplicator(310), ---  -0.757202148438
            im_multiplicator => im_multiplicator(310), --- j-0.653198242188
            data_re_out => mul_re_out(310),
            data_im_out => mul_im_out(310)
        );

 
    UMUL_311 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(311),
            data_im_in => first_stage_im_out(311),
            re_multiplicator => re_multiplicator(311), ---  -0.824584960938
            im_multiplicator => im_multiplicator(311), --- j-0.565734863281
            data_re_out => mul_re_out(311),
            data_im_out => mul_im_out(311)
        );

 
    UMUL_312 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(312),
            data_im_in => first_stage_im_out(312),
            re_multiplicator => re_multiplicator(312), ---  -0.881896972656
            im_multiplicator => im_multiplicator(312), --- j-0.471374511719
            data_re_out => mul_re_out(312),
            data_im_out => mul_im_out(312)
        );

 
    UMUL_313 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(313),
            data_im_in => first_stage_im_out(313),
            re_multiplicator => re_multiplicator(313), ---  -0.928527832031
            im_multiplicator => im_multiplicator(313), --- j-0.371337890625
            data_re_out => mul_re_out(313),
            data_im_out => mul_im_out(313)
        );

 
    UMUL_314 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(314),
            data_im_in => first_stage_im_out(314),
            re_multiplicator => re_multiplicator(314), ---  -0.963806152344
            im_multiplicator => im_multiplicator(314), --- j-0.266723632812
            data_re_out => mul_re_out(314),
            data_im_out => mul_im_out(314)
        );

 
    UMUL_315 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(315),
            data_im_in => first_stage_im_out(315),
            re_multiplicator => re_multiplicator(315), ---  -0.9873046875
            im_multiplicator => im_multiplicator(315), --- j-0.158874511719
            data_re_out => mul_re_out(315),
            data_im_out => mul_im_out(315)
        );

 
    UMUL_316 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(316),
            data_im_in => first_stage_im_out(316),
            re_multiplicator => re_multiplicator(316), ---  -0.998779296875
            im_multiplicator => im_multiplicator(316), --- j-0.049072265625
            data_re_out => mul_re_out(316),
            data_im_out => mul_im_out(316)
        );

 
    UMUL_317 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(317),
            data_im_in => first_stage_im_out(317),
            re_multiplicator => re_multiplicator(317), ---  -0.998107910156
            im_multiplicator => im_multiplicator(317), --- j0.0613403320312
            data_re_out => mul_re_out(317),
            data_im_out => mul_im_out(317)
        );

 
    UMUL_318 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(318),
            data_im_in => first_stage_im_out(318),
            re_multiplicator => re_multiplicator(318), ---  -0.985290527344
            im_multiplicator => im_multiplicator(318), --- j0.170959472656
            data_re_out => mul_re_out(318),
            data_im_out => mul_im_out(318)
        );

 
    UMUL_319 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(319),
            data_im_in => first_stage_im_out(319),
            re_multiplicator => re_multiplicator(319), ---  -0.96044921875
            im_multiplicator => im_multiplicator(319), --- j0.278503417969
            data_re_out => mul_re_out(319),
            data_im_out => mul_im_out(319)
        );

 
    UMUL_320 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(320),
            data_im_in => first_stage_im_out(320),
            data_re_out => mul_re_out(320),
            data_im_out => mul_im_out(320)
        );

 
    UMUL_321 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(321),
            data_im_in => first_stage_im_out(321),
            re_multiplicator => re_multiplicator(321), ---  0.992492675781
            im_multiplicator => im_multiplicator(321), --- j-0.122436523438
            data_re_out => mul_re_out(321),
            data_im_out => mul_im_out(321)
        );

 
    UMUL_322 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(322),
            data_im_in => first_stage_im_out(322),
            re_multiplicator => re_multiplicator(322), ---  0.970031738281
            im_multiplicator => im_multiplicator(322), --- j-0.242980957031
            data_re_out => mul_re_out(322),
            data_im_out => mul_im_out(322)
        );

 
    UMUL_323 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(323),
            data_im_in => first_stage_im_out(323),
            re_multiplicator => re_multiplicator(323), ---  0.932983398438
            im_multiplicator => im_multiplicator(323), --- j-0.359924316406
            data_re_out => mul_re_out(323),
            data_im_out => mul_im_out(323)
        );

 
    UMUL_324 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(324),
            data_im_in => first_stage_im_out(324),
            re_multiplicator => re_multiplicator(324), ---  0.881896972656
            im_multiplicator => im_multiplicator(324), --- j-0.471374511719
            data_re_out => mul_re_out(324),
            data_im_out => mul_im_out(324)
        );

 
    UMUL_325 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(325),
            data_im_in => first_stage_im_out(325),
            re_multiplicator => re_multiplicator(325), ---  0.817565917969
            im_multiplicator => im_multiplicator(325), --- j-0.575805664062
            data_re_out => mul_re_out(325),
            data_im_out => mul_im_out(325)
        );

 
    UMUL_326 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(326),
            data_im_in => first_stage_im_out(326),
            re_multiplicator => re_multiplicator(326), ---  0.740966796875
            im_multiplicator => im_multiplicator(326), --- j-0.671569824219
            data_re_out => mul_re_out(326),
            data_im_out => mul_im_out(326)
        );

 
    UMUL_327 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(327),
            data_im_in => first_stage_im_out(327),
            re_multiplicator => re_multiplicator(327), ---  0.653198242188
            im_multiplicator => im_multiplicator(327), --- j-0.757202148438
            data_re_out => mul_re_out(327),
            data_im_out => mul_im_out(327)
        );

 
    UMUL_328 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(328),
            data_im_in => first_stage_im_out(328),
            re_multiplicator => re_multiplicator(328), ---  0.555541992188
            im_multiplicator => im_multiplicator(328), --- j-0.831481933594
            data_re_out => mul_re_out(328),
            data_im_out => mul_im_out(328)
        );

 
    UMUL_329 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(329),
            data_im_in => first_stage_im_out(329),
            re_multiplicator => re_multiplicator(329), ---  0.449584960938
            im_multiplicator => im_multiplicator(329), --- j-0.893249511719
            data_re_out => mul_re_out(329),
            data_im_out => mul_im_out(329)
        );

 
    UMUL_330 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(330),
            data_im_in => first_stage_im_out(330),
            re_multiplicator => re_multiplicator(330), ---  0.3369140625
            im_multiplicator => im_multiplicator(330), --- j-0.941528320312
            data_re_out => mul_re_out(330),
            data_im_out => mul_im_out(330)
        );

 
    UMUL_331 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(331),
            data_im_in => first_stage_im_out(331),
            re_multiplicator => re_multiplicator(331), ---  0.219116210938
            im_multiplicator => im_multiplicator(331), --- j-0.975708007812
            data_re_out => mul_re_out(331),
            data_im_out => mul_im_out(331)
        );

 
    UMUL_332 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(332),
            data_im_in => first_stage_im_out(332),
            re_multiplicator => re_multiplicator(332), ---  0.0980224609375
            im_multiplicator => im_multiplicator(332), --- j-0.995178222656
            data_re_out => mul_re_out(332),
            data_im_out => mul_im_out(332)
        );

 
    UMUL_333 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(333),
            data_im_in => first_stage_im_out(333),
            re_multiplicator => re_multiplicator(333), ---  -0.0245361328125
            im_multiplicator => im_multiplicator(333), --- j-0.999694824219
            data_re_out => mul_re_out(333),
            data_im_out => mul_im_out(333)
        );

 
    UMUL_334 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(334),
            data_im_in => first_stage_im_out(334),
            re_multiplicator => re_multiplicator(334), ---  -0.146728515625
            im_multiplicator => im_multiplicator(334), --- j-0.989196777344
            data_re_out => mul_re_out(334),
            data_im_out => mul_im_out(334)
        );

 
    UMUL_335 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(335),
            data_im_in => first_stage_im_out(335),
            re_multiplicator => re_multiplicator(335), ---  -0.266723632812
            im_multiplicator => im_multiplicator(335), --- j-0.963806152344
            data_re_out => mul_re_out(335),
            data_im_out => mul_im_out(335)
        );

 
    UMUL_336 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(336),
            data_im_in => first_stage_im_out(336),
            re_multiplicator => re_multiplicator(336), ---  -0.382690429688
            im_multiplicator => im_multiplicator(336), --- j-0.923889160156
            data_re_out => mul_re_out(336),
            data_im_out => mul_im_out(336)
        );

 
    UMUL_337 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(337),
            data_im_in => first_stage_im_out(337),
            re_multiplicator => re_multiplicator(337), ---  -0.492919921875
            im_multiplicator => im_multiplicator(337), --- j-0.8701171875
            data_re_out => mul_re_out(337),
            data_im_out => mul_im_out(337)
        );

 
    UMUL_338 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(338),
            data_im_in => first_stage_im_out(338),
            re_multiplicator => re_multiplicator(338), ---  -0.595703125
            im_multiplicator => im_multiplicator(338), --- j-0.80322265625
            data_re_out => mul_re_out(338),
            data_im_out => mul_im_out(338)
        );

 
    UMUL_339 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(339),
            data_im_in => first_stage_im_out(339),
            re_multiplicator => re_multiplicator(339), ---  -0.689514160156
            im_multiplicator => im_multiplicator(339), --- j-0.724243164062
            data_re_out => mul_re_out(339),
            data_im_out => mul_im_out(339)
        );

 
    UMUL_340 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(340),
            data_im_in => first_stage_im_out(340),
            re_multiplicator => re_multiplicator(340), ---  -0.773010253906
            im_multiplicator => im_multiplicator(340), --- j-0.634399414062
            data_re_out => mul_re_out(340),
            data_im_out => mul_im_out(340)
        );

 
    UMUL_341 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(341),
            data_im_in => first_stage_im_out(341),
            re_multiplicator => re_multiplicator(341), ---  -0.844848632812
            im_multiplicator => im_multiplicator(341), --- j-0.534973144531
            data_re_out => mul_re_out(341),
            data_im_out => mul_im_out(341)
        );

 
    UMUL_342 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(342),
            data_im_in => first_stage_im_out(342),
            re_multiplicator => re_multiplicator(342), ---  -0.903991699219
            im_multiplicator => im_multiplicator(342), --- j-0.427551269531
            data_re_out => mul_re_out(342),
            data_im_out => mul_im_out(342)
        );

 
    UMUL_343 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(343),
            data_im_in => first_stage_im_out(343),
            re_multiplicator => re_multiplicator(343), ---  -0.949523925781
            im_multiplicator => im_multiplicator(343), --- j-0.313659667969
            data_re_out => mul_re_out(343),
            data_im_out => mul_im_out(343)
        );

 
    UMUL_344 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(344),
            data_im_in => first_stage_im_out(344),
            re_multiplicator => re_multiplicator(344), ---  -0.980773925781
            im_multiplicator => im_multiplicator(344), --- j-0.195068359375
            data_re_out => mul_re_out(344),
            data_im_out => mul_im_out(344)
        );

 
    UMUL_345 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(345),
            data_im_in => first_stage_im_out(345),
            re_multiplicator => re_multiplicator(345), ---  -0.997314453125
            im_multiplicator => im_multiplicator(345), --- j-0.0735473632812
            data_re_out => mul_re_out(345),
            data_im_out => mul_im_out(345)
        );

 
    UMUL_346 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(346),
            data_im_in => first_stage_im_out(346),
            re_multiplicator => re_multiplicator(346), ---  -0.998779296875
            im_multiplicator => im_multiplicator(346), --- j0.049072265625
            data_re_out => mul_re_out(346),
            data_im_out => mul_im_out(346)
        );

 
    UMUL_347 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(347),
            data_im_in => first_stage_im_out(347),
            re_multiplicator => re_multiplicator(347), ---  -0.985290527344
            im_multiplicator => im_multiplicator(347), --- j0.170959472656
            data_re_out => mul_re_out(347),
            data_im_out => mul_im_out(347)
        );

 
    UMUL_348 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(348),
            data_im_in => first_stage_im_out(348),
            re_multiplicator => re_multiplicator(348), ---  -0.956970214844
            im_multiplicator => im_multiplicator(348), --- j0.290283203125
            data_re_out => mul_re_out(348),
            data_im_out => mul_im_out(348)
        );

 
    UMUL_349 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(349),
            data_im_in => first_stage_im_out(349),
            re_multiplicator => re_multiplicator(349), ---  -0.914184570312
            im_multiplicator => im_multiplicator(349), --- j0.405212402344
            data_re_out => mul_re_out(349),
            data_im_out => mul_im_out(349)
        );

 
    UMUL_350 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(350),
            data_im_in => first_stage_im_out(350),
            re_multiplicator => re_multiplicator(350), ---  -0.857727050781
            im_multiplicator => im_multiplicator(350), --- j0.514099121094
            data_re_out => mul_re_out(350),
            data_im_out => mul_im_out(350)
        );

 
    UMUL_351 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(351),
            data_im_in => first_stage_im_out(351),
            re_multiplicator => re_multiplicator(351), ---  -0.788330078125
            im_multiplicator => im_multiplicator(351), --- j0.615234375
            data_re_out => mul_re_out(351),
            data_im_out => mul_im_out(351)
        );

 
    UMUL_352 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(352),
            data_im_in => first_stage_im_out(352),
            data_re_out => mul_re_out(352),
            data_im_out => mul_im_out(352)
        );

 
    UMUL_353 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(353),
            data_im_in => first_stage_im_out(353),
            re_multiplicator => re_multiplicator(353), ---  0.990905761719
            im_multiplicator => im_multiplicator(353), --- j-0.134582519531
            data_re_out => mul_re_out(353),
            data_im_out => mul_im_out(353)
        );

 
    UMUL_354 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(354),
            data_im_in => first_stage_im_out(354),
            re_multiplicator => re_multiplicator(354), ---  0.963806152344
            im_multiplicator => im_multiplicator(354), --- j-0.266723632812
            data_re_out => mul_re_out(354),
            data_im_out => mul_im_out(354)
        );

 
    UMUL_355 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(355),
            data_im_in => first_stage_im_out(355),
            re_multiplicator => re_multiplicator(355), ---  0.919128417969
            im_multiplicator => im_multiplicator(355), --- j-0.393981933594
            data_re_out => mul_re_out(355),
            data_im_out => mul_im_out(355)
        );

 
    UMUL_356 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(356),
            data_im_in => first_stage_im_out(356),
            re_multiplicator => re_multiplicator(356), ---  0.857727050781
            im_multiplicator => im_multiplicator(356), --- j-0.514099121094
            data_re_out => mul_re_out(356),
            data_im_out => mul_im_out(356)
        );

 
    UMUL_357 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(357),
            data_im_in => first_stage_im_out(357),
            re_multiplicator => re_multiplicator(357), ---  0.78076171875
            im_multiplicator => im_multiplicator(357), --- j-0.624877929688
            data_re_out => mul_re_out(357),
            data_im_out => mul_im_out(357)
        );

 
    UMUL_358 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(358),
            data_im_in => first_stage_im_out(358),
            re_multiplicator => re_multiplicator(358), ---  0.689514160156
            im_multiplicator => im_multiplicator(358), --- j-0.724243164062
            data_re_out => mul_re_out(358),
            data_im_out => mul_im_out(358)
        );

 
    UMUL_359 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(359),
            data_im_in => first_stage_im_out(359),
            re_multiplicator => re_multiplicator(359), ---  0.585815429688
            im_multiplicator => im_multiplicator(359), --- j-0.810485839844
            data_re_out => mul_re_out(359),
            data_im_out => mul_im_out(359)
        );

 
    UMUL_360 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(360),
            data_im_in => first_stage_im_out(360),
            re_multiplicator => re_multiplicator(360), ---  0.471374511719
            im_multiplicator => im_multiplicator(360), --- j-0.881896972656
            data_re_out => mul_re_out(360),
            data_im_out => mul_im_out(360)
        );

 
    UMUL_361 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(361),
            data_im_in => first_stage_im_out(361),
            re_multiplicator => re_multiplicator(361), ---  0.348388671875
            im_multiplicator => im_multiplicator(361), --- j-0.937316894531
            data_re_out => mul_re_out(361),
            data_im_out => mul_im_out(361)
        );

 
    UMUL_362 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(362),
            data_im_in => first_stage_im_out(362),
            re_multiplicator => re_multiplicator(362), ---  0.219116210938
            im_multiplicator => im_multiplicator(362), --- j-0.975708007812
            data_re_out => mul_re_out(362),
            data_im_out => mul_im_out(362)
        );

 
    UMUL_363 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(363),
            data_im_in => first_stage_im_out(363),
            re_multiplicator => re_multiplicator(363), ---  0.0858154296875
            im_multiplicator => im_multiplicator(363), --- j-0.996337890625
            data_re_out => mul_re_out(363),
            data_im_out => mul_im_out(363)
        );

 
    UMUL_364 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(364),
            data_im_in => first_stage_im_out(364),
            re_multiplicator => re_multiplicator(364), ---  -0.049072265625
            im_multiplicator => im_multiplicator(364), --- j-0.998779296875
            data_re_out => mul_re_out(364),
            data_im_out => mul_im_out(364)
        );

 
    UMUL_365 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(365),
            data_im_in => first_stage_im_out(365),
            re_multiplicator => re_multiplicator(365), ---  -0.183044433594
            im_multiplicator => im_multiplicator(365), --- j-0.983093261719
            data_re_out => mul_re_out(365),
            data_im_out => mul_im_out(365)
        );

 
    UMUL_366 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(366),
            data_im_in => first_stage_im_out(366),
            re_multiplicator => re_multiplicator(366), ---  -0.313659667969
            im_multiplicator => im_multiplicator(366), --- j-0.949523925781
            data_re_out => mul_re_out(366),
            data_im_out => mul_im_out(366)
        );

 
    UMUL_367 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(367),
            data_im_in => first_stage_im_out(367),
            re_multiplicator => re_multiplicator(367), ---  -0.438598632812
            im_multiplicator => im_multiplicator(367), --- j-0.898681640625
            data_re_out => mul_re_out(367),
            data_im_out => mul_im_out(367)
        );

 
    UMUL_368 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(368),
            data_im_in => first_stage_im_out(368),
            re_multiplicator => re_multiplicator(368), ---  -0.555541992188
            im_multiplicator => im_multiplicator(368), --- j-0.831481933594
            data_re_out => mul_re_out(368),
            data_im_out => mul_im_out(368)
        );

 
    UMUL_369 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(369),
            data_im_in => first_stage_im_out(369),
            re_multiplicator => re_multiplicator(369), ---  -0.662414550781
            im_multiplicator => im_multiplicator(369), --- j-0.749145507812
            data_re_out => mul_re_out(369),
            data_im_out => mul_im_out(369)
        );

 
    UMUL_370 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(370),
            data_im_in => first_stage_im_out(370),
            re_multiplicator => re_multiplicator(370), ---  -0.757202148438
            im_multiplicator => im_multiplicator(370), --- j-0.653198242188
            data_re_out => mul_re_out(370),
            data_im_out => mul_im_out(370)
        );

 
    UMUL_371 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(371),
            data_im_in => first_stage_im_out(371),
            re_multiplicator => re_multiplicator(371), ---  -0.838195800781
            im_multiplicator => im_multiplicator(371), --- j-0.545349121094
            data_re_out => mul_re_out(371),
            data_im_out => mul_im_out(371)
        );

 
    UMUL_372 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(372),
            data_im_in => first_stage_im_out(372),
            re_multiplicator => re_multiplicator(372), ---  -0.903991699219
            im_multiplicator => im_multiplicator(372), --- j-0.427551269531
            data_re_out => mul_re_out(372),
            data_im_out => mul_im_out(372)
        );

 
    UMUL_373 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(373),
            data_im_in => first_stage_im_out(373),
            re_multiplicator => re_multiplicator(373), ---  -0.953308105469
            im_multiplicator => im_multiplicator(373), --- j-0.302001953125
            data_re_out => mul_re_out(373),
            data_im_out => mul_im_out(373)
        );

 
    UMUL_374 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(374),
            data_im_in => first_stage_im_out(374),
            re_multiplicator => re_multiplicator(374), ---  -0.985290527344
            im_multiplicator => im_multiplicator(374), --- j-0.170959472656
            data_re_out => mul_re_out(374),
            data_im_out => mul_im_out(374)
        );

 
    UMUL_375 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(375),
            data_im_in => first_stage_im_out(375),
            re_multiplicator => re_multiplicator(375), ---  -0.999328613281
            im_multiplicator => im_multiplicator(375), --- j-0.0368041992188
            data_re_out => mul_re_out(375),
            data_im_out => mul_im_out(375)
        );

 
    UMUL_376 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(376),
            data_im_in => first_stage_im_out(376),
            re_multiplicator => re_multiplicator(376), ---  -0.995178222656
            im_multiplicator => im_multiplicator(376), --- j0.0980224609375
            data_re_out => mul_re_out(376),
            data_im_out => mul_im_out(376)
        );

 
    UMUL_377 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(377),
            data_im_in => first_stage_im_out(377),
            re_multiplicator => re_multiplicator(377), ---  -0.972961425781
            im_multiplicator => im_multiplicator(377), --- j0.231079101562
            data_re_out => mul_re_out(377),
            data_im_out => mul_im_out(377)
        );

 
    UMUL_378 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(378),
            data_im_in => first_stage_im_out(378),
            re_multiplicator => re_multiplicator(378), ---  -0.932983398438
            im_multiplicator => im_multiplicator(378), --- j0.359924316406
            data_re_out => mul_re_out(378),
            data_im_out => mul_im_out(378)
        );

 
    UMUL_379 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(379),
            data_im_in => first_stage_im_out(379),
            re_multiplicator => re_multiplicator(379), ---  -0.876098632812
            im_multiplicator => im_multiplicator(379), --- j0.482177734375
            data_re_out => mul_re_out(379),
            data_im_out => mul_im_out(379)
        );

 
    UMUL_380 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(380),
            data_im_in => first_stage_im_out(380),
            re_multiplicator => re_multiplicator(380), ---  -0.80322265625
            im_multiplicator => im_multiplicator(380), --- j0.595703125
            data_re_out => mul_re_out(380),
            data_im_out => mul_im_out(380)
        );

 
    UMUL_381 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(381),
            data_im_in => first_stage_im_out(381),
            re_multiplicator => re_multiplicator(381), ---  -0.715759277344
            im_multiplicator => im_multiplicator(381), --- j0.698364257812
            data_re_out => mul_re_out(381),
            data_im_out => mul_im_out(381)
        );

 
    UMUL_382 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(382),
            data_im_in => first_stage_im_out(382),
            re_multiplicator => re_multiplicator(382), ---  -0.615234375
            im_multiplicator => im_multiplicator(382), --- j0.788330078125
            data_re_out => mul_re_out(382),
            data_im_out => mul_im_out(382)
        );

 
    UMUL_383 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(383),
            data_im_in => first_stage_im_out(383),
            re_multiplicator => re_multiplicator(383), ---  -0.503540039062
            im_multiplicator => im_multiplicator(383), --- j0.863952636719
            data_re_out => mul_re_out(383),
            data_im_out => mul_im_out(383)
        );

 
    UMUL_384 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(384),
            data_im_in => first_stage_im_out(384),
            data_re_out => mul_re_out(384),
            data_im_out => mul_im_out(384)
        );

 
    UMUL_385 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(385),
            data_im_in => first_stage_im_out(385),
            re_multiplicator => re_multiplicator(385), ---  0.989196777344
            im_multiplicator => im_multiplicator(385), --- j-0.146728515625
            data_re_out => mul_re_out(385),
            data_im_out => mul_im_out(385)
        );

 
    UMUL_386 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(386),
            data_im_in => first_stage_im_out(386),
            re_multiplicator => re_multiplicator(386), ---  0.956970214844
            im_multiplicator => im_multiplicator(386), --- j-0.290283203125
            data_re_out => mul_re_out(386),
            data_im_out => mul_im_out(386)
        );

 
    UMUL_387 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(387),
            data_im_in => first_stage_im_out(387),
            re_multiplicator => re_multiplicator(387), ---  0.903991699219
            im_multiplicator => im_multiplicator(387), --- j-0.427551269531
            data_re_out => mul_re_out(387),
            data_im_out => mul_im_out(387)
        );

 
    UMUL_388 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(388),
            data_im_in => first_stage_im_out(388),
            re_multiplicator => re_multiplicator(388), ---  0.831481933594
            im_multiplicator => im_multiplicator(388), --- j-0.555541992188
            data_re_out => mul_re_out(388),
            data_im_out => mul_im_out(388)
        );

 
    UMUL_389 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(389),
            data_im_in => first_stage_im_out(389),
            re_multiplicator => re_multiplicator(389), ---  0.740966796875
            im_multiplicator => im_multiplicator(389), --- j-0.671569824219
            data_re_out => mul_re_out(389),
            data_im_out => mul_im_out(389)
        );

 
    UMUL_390 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(390),
            data_im_in => first_stage_im_out(390),
            re_multiplicator => re_multiplicator(390), ---  0.634399414062
            im_multiplicator => im_multiplicator(390), --- j-0.773010253906
            data_re_out => mul_re_out(390),
            data_im_out => mul_im_out(390)
        );

 
    UMUL_391 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(391),
            data_im_in => first_stage_im_out(391),
            re_multiplicator => re_multiplicator(391), ---  0.514099121094
            im_multiplicator => im_multiplicator(391), --- j-0.857727050781
            data_re_out => mul_re_out(391),
            data_im_out => mul_im_out(391)
        );

 
    UMUL_392 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(392),
            data_im_in => first_stage_im_out(392),
            re_multiplicator => re_multiplicator(392), ---  0.382690429688
            im_multiplicator => im_multiplicator(392), --- j-0.923889160156
            data_re_out => mul_re_out(392),
            data_im_out => mul_im_out(392)
        );

 
    UMUL_393 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(393),
            data_im_in => first_stage_im_out(393),
            re_multiplicator => re_multiplicator(393), ---  0.242980957031
            im_multiplicator => im_multiplicator(393), --- j-0.970031738281
            data_re_out => mul_re_out(393),
            data_im_out => mul_im_out(393)
        );

 
    UMUL_394 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(394),
            data_im_in => first_stage_im_out(394),
            re_multiplicator => re_multiplicator(394), ---  0.0980224609375
            im_multiplicator => im_multiplicator(394), --- j-0.995178222656
            data_re_out => mul_re_out(394),
            data_im_out => mul_im_out(394)
        );

 
    UMUL_395 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(395),
            data_im_in => first_stage_im_out(395),
            re_multiplicator => re_multiplicator(395), ---  -0.049072265625
            im_multiplicator => im_multiplicator(395), --- j-0.998779296875
            data_re_out => mul_re_out(395),
            data_im_out => mul_im_out(395)
        );

 
    UMUL_396 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(396),
            data_im_in => first_stage_im_out(396),
            re_multiplicator => re_multiplicator(396), ---  -0.195068359375
            im_multiplicator => im_multiplicator(396), --- j-0.980773925781
            data_re_out => mul_re_out(396),
            data_im_out => mul_im_out(396)
        );

 
    UMUL_397 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(397),
            data_im_in => first_stage_im_out(397),
            re_multiplicator => re_multiplicator(397), ---  -0.3369140625
            im_multiplicator => im_multiplicator(397), --- j-0.941528320312
            data_re_out => mul_re_out(397),
            data_im_out => mul_im_out(397)
        );

 
    UMUL_398 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(398),
            data_im_in => first_stage_im_out(398),
            re_multiplicator => re_multiplicator(398), ---  -0.471374511719
            im_multiplicator => im_multiplicator(398), --- j-0.881896972656
            data_re_out => mul_re_out(398),
            data_im_out => mul_im_out(398)
        );

 
    UMUL_399 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(399),
            data_im_in => first_stage_im_out(399),
            re_multiplicator => re_multiplicator(399), ---  -0.595703125
            im_multiplicator => im_multiplicator(399), --- j-0.80322265625
            data_re_out => mul_re_out(399),
            data_im_out => mul_im_out(399)
        );

 
    UMUL_400 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(400),
            data_im_in => first_stage_im_out(400),
            re_multiplicator => re_multiplicator(400), ---  -0.707092285156
            im_multiplicator => im_multiplicator(400), --- j-0.707092285156
            data_re_out => mul_re_out(400),
            data_im_out => mul_im_out(400)
        );

 
    UMUL_401 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(401),
            data_im_in => first_stage_im_out(401),
            re_multiplicator => re_multiplicator(401), ---  -0.80322265625
            im_multiplicator => im_multiplicator(401), --- j-0.595703125
            data_re_out => mul_re_out(401),
            data_im_out => mul_im_out(401)
        );

 
    UMUL_402 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(402),
            data_im_in => first_stage_im_out(402),
            re_multiplicator => re_multiplicator(402), ---  -0.881896972656
            im_multiplicator => im_multiplicator(402), --- j-0.471374511719
            data_re_out => mul_re_out(402),
            data_im_out => mul_im_out(402)
        );

 
    UMUL_403 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(403),
            data_im_in => first_stage_im_out(403),
            re_multiplicator => re_multiplicator(403), ---  -0.941528320312
            im_multiplicator => im_multiplicator(403), --- j-0.3369140625
            data_re_out => mul_re_out(403),
            data_im_out => mul_im_out(403)
        );

 
    UMUL_404 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(404),
            data_im_in => first_stage_im_out(404),
            re_multiplicator => re_multiplicator(404), ---  -0.980773925781
            im_multiplicator => im_multiplicator(404), --- j-0.195068359375
            data_re_out => mul_re_out(404),
            data_im_out => mul_im_out(404)
        );

 
    UMUL_405 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(405),
            data_im_in => first_stage_im_out(405),
            re_multiplicator => re_multiplicator(405), ---  -0.998779296875
            im_multiplicator => im_multiplicator(405), --- j-0.049072265625
            data_re_out => mul_re_out(405),
            data_im_out => mul_im_out(405)
        );

 
    UMUL_406 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(406),
            data_im_in => first_stage_im_out(406),
            re_multiplicator => re_multiplicator(406), ---  -0.995178222656
            im_multiplicator => im_multiplicator(406), --- j0.0980224609375
            data_re_out => mul_re_out(406),
            data_im_out => mul_im_out(406)
        );

 
    UMUL_407 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(407),
            data_im_in => first_stage_im_out(407),
            re_multiplicator => re_multiplicator(407), ---  -0.970031738281
            im_multiplicator => im_multiplicator(407), --- j0.242980957031
            data_re_out => mul_re_out(407),
            data_im_out => mul_im_out(407)
        );

 
    UMUL_408 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(408),
            data_im_in => first_stage_im_out(408),
            re_multiplicator => re_multiplicator(408), ---  -0.923889160156
            im_multiplicator => im_multiplicator(408), --- j0.382690429688
            data_re_out => mul_re_out(408),
            data_im_out => mul_im_out(408)
        );

 
    UMUL_409 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(409),
            data_im_in => first_stage_im_out(409),
            re_multiplicator => re_multiplicator(409), ---  -0.857727050781
            im_multiplicator => im_multiplicator(409), --- j0.514099121094
            data_re_out => mul_re_out(409),
            data_im_out => mul_im_out(409)
        );

 
    UMUL_410 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(410),
            data_im_in => first_stage_im_out(410),
            re_multiplicator => re_multiplicator(410), ---  -0.773010253906
            im_multiplicator => im_multiplicator(410), --- j0.634399414062
            data_re_out => mul_re_out(410),
            data_im_out => mul_im_out(410)
        );

 
    UMUL_411 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(411),
            data_im_in => first_stage_im_out(411),
            re_multiplicator => re_multiplicator(411), ---  -0.671569824219
            im_multiplicator => im_multiplicator(411), --- j0.740966796875
            data_re_out => mul_re_out(411),
            data_im_out => mul_im_out(411)
        );

 
    UMUL_412 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(412),
            data_im_in => first_stage_im_out(412),
            re_multiplicator => re_multiplicator(412), ---  -0.555541992188
            im_multiplicator => im_multiplicator(412), --- j0.831481933594
            data_re_out => mul_re_out(412),
            data_im_out => mul_im_out(412)
        );

 
    UMUL_413 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(413),
            data_im_in => first_stage_im_out(413),
            re_multiplicator => re_multiplicator(413), ---  -0.427551269531
            im_multiplicator => im_multiplicator(413), --- j0.903991699219
            data_re_out => mul_re_out(413),
            data_im_out => mul_im_out(413)
        );

 
    UMUL_414 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(414),
            data_im_in => first_stage_im_out(414),
            re_multiplicator => re_multiplicator(414), ---  -0.290283203125
            im_multiplicator => im_multiplicator(414), --- j0.956970214844
            data_re_out => mul_re_out(414),
            data_im_out => mul_im_out(414)
        );

 
    UMUL_415 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(415),
            data_im_in => first_stage_im_out(415),
            re_multiplicator => re_multiplicator(415), ---  -0.146728515625
            im_multiplicator => im_multiplicator(415), --- j0.989196777344
            data_re_out => mul_re_out(415),
            data_im_out => mul_im_out(415)
        );

 
    UMUL_416 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(416),
            data_im_in => first_stage_im_out(416),
            data_re_out => mul_re_out(416),
            data_im_out => mul_im_out(416)
        );

 
    UMUL_417 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(417),
            data_im_in => first_stage_im_out(417),
            re_multiplicator => re_multiplicator(417), ---  0.9873046875
            im_multiplicator => im_multiplicator(417), --- j-0.158874511719
            data_re_out => mul_re_out(417),
            data_im_out => mul_im_out(417)
        );

 
    UMUL_418 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(418),
            data_im_in => first_stage_im_out(418),
            re_multiplicator => re_multiplicator(418), ---  0.949523925781
            im_multiplicator => im_multiplicator(418), --- j-0.313659667969
            data_re_out => mul_re_out(418),
            data_im_out => mul_im_out(418)
        );

 
    UMUL_419 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(419),
            data_im_in => first_stage_im_out(419),
            re_multiplicator => re_multiplicator(419), ---  0.887634277344
            im_multiplicator => im_multiplicator(419), --- j-0.460510253906
            data_re_out => mul_re_out(419),
            data_im_out => mul_im_out(419)
        );

 
    UMUL_420 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(420),
            data_im_in => first_stage_im_out(420),
            re_multiplicator => re_multiplicator(420), ---  0.80322265625
            im_multiplicator => im_multiplicator(420), --- j-0.595703125
            data_re_out => mul_re_out(420),
            data_im_out => mul_im_out(420)
        );

 
    UMUL_421 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(421),
            data_im_in => first_stage_im_out(421),
            re_multiplicator => re_multiplicator(421), ---  0.698364257812
            im_multiplicator => im_multiplicator(421), --- j-0.715759277344
            data_re_out => mul_re_out(421),
            data_im_out => mul_im_out(421)
        );

 
    UMUL_422 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(422),
            data_im_in => first_stage_im_out(422),
            re_multiplicator => re_multiplicator(422), ---  0.575805664062
            im_multiplicator => im_multiplicator(422), --- j-0.817565917969
            data_re_out => mul_re_out(422),
            data_im_out => mul_im_out(422)
        );

 
    UMUL_423 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(423),
            data_im_in => first_stage_im_out(423),
            re_multiplicator => re_multiplicator(423), ---  0.438598632812
            im_multiplicator => im_multiplicator(423), --- j-0.898681640625
            data_re_out => mul_re_out(423),
            data_im_out => mul_im_out(423)
        );

 
    UMUL_424 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(424),
            data_im_in => first_stage_im_out(424),
            re_multiplicator => re_multiplicator(424), ---  0.290283203125
            im_multiplicator => im_multiplicator(424), --- j-0.956970214844
            data_re_out => mul_re_out(424),
            data_im_out => mul_im_out(424)
        );

 
    UMUL_425 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(425),
            data_im_in => first_stage_im_out(425),
            re_multiplicator => re_multiplicator(425), ---  0.134582519531
            im_multiplicator => im_multiplicator(425), --- j-0.990905761719
            data_re_out => mul_re_out(425),
            data_im_out => mul_im_out(425)
        );

 
    UMUL_426 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(426),
            data_im_in => first_stage_im_out(426),
            re_multiplicator => re_multiplicator(426), ---  -0.0245361328125
            im_multiplicator => im_multiplicator(426), --- j-0.999694824219
            data_re_out => mul_re_out(426),
            data_im_out => mul_im_out(426)
        );

 
    UMUL_427 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(427),
            data_im_in => first_stage_im_out(427),
            re_multiplicator => re_multiplicator(427), ---  -0.183044433594
            im_multiplicator => im_multiplicator(427), --- j-0.983093261719
            data_re_out => mul_re_out(427),
            data_im_out => mul_im_out(427)
        );

 
    UMUL_428 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(428),
            data_im_in => first_stage_im_out(428),
            re_multiplicator => re_multiplicator(428), ---  -0.3369140625
            im_multiplicator => im_multiplicator(428), --- j-0.941528320312
            data_re_out => mul_re_out(428),
            data_im_out => mul_im_out(428)
        );

 
    UMUL_429 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(429),
            data_im_in => first_stage_im_out(429),
            re_multiplicator => re_multiplicator(429), ---  -0.482177734375
            im_multiplicator => im_multiplicator(429), --- j-0.876098632812
            data_re_out => mul_re_out(429),
            data_im_out => mul_im_out(429)
        );

 
    UMUL_430 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(430),
            data_im_in => first_stage_im_out(430),
            re_multiplicator => re_multiplicator(430), ---  -0.615234375
            im_multiplicator => im_multiplicator(430), --- j-0.788330078125
            data_re_out => mul_re_out(430),
            data_im_out => mul_im_out(430)
        );

 
    UMUL_431 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(431),
            data_im_in => first_stage_im_out(431),
            re_multiplicator => re_multiplicator(431), ---  -0.732666015625
            im_multiplicator => im_multiplicator(431), --- j-0.680603027344
            data_re_out => mul_re_out(431),
            data_im_out => mul_im_out(431)
        );

 
    UMUL_432 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(432),
            data_im_in => first_stage_im_out(432),
            re_multiplicator => re_multiplicator(432), ---  -0.831481933594
            im_multiplicator => im_multiplicator(432), --- j-0.555541992188
            data_re_out => mul_re_out(432),
            data_im_out => mul_im_out(432)
        );

 
    UMUL_433 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(433),
            data_im_in => first_stage_im_out(433),
            re_multiplicator => re_multiplicator(433), ---  -0.9091796875
            im_multiplicator => im_multiplicator(433), --- j-0.416442871094
            data_re_out => mul_re_out(433),
            data_im_out => mul_im_out(433)
        );

 
    UMUL_434 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(434),
            data_im_in => first_stage_im_out(434),
            re_multiplicator => re_multiplicator(434), ---  -0.963806152344
            im_multiplicator => im_multiplicator(434), --- j-0.266723632812
            data_re_out => mul_re_out(434),
            data_im_out => mul_im_out(434)
        );

 
    UMUL_435 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(435),
            data_im_in => first_stage_im_out(435),
            re_multiplicator => re_multiplicator(435), ---  -0.993896484375
            im_multiplicator => im_multiplicator(435), --- j-0.110229492188
            data_re_out => mul_re_out(435),
            data_im_out => mul_im_out(435)
        );

 
    UMUL_436 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(436),
            data_im_in => first_stage_im_out(436),
            re_multiplicator => re_multiplicator(436), ---  -0.998779296875
            im_multiplicator => im_multiplicator(436), --- j0.049072265625
            data_re_out => mul_re_out(436),
            data_im_out => mul_im_out(436)
        );

 
    UMUL_437 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(437),
            data_im_in => first_stage_im_out(437),
            re_multiplicator => re_multiplicator(437), ---  -0.978332519531
            im_multiplicator => im_multiplicator(437), --- j0.207092285156
            data_re_out => mul_re_out(437),
            data_im_out => mul_im_out(437)
        );

 
    UMUL_438 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(438),
            data_im_in => first_stage_im_out(438),
            re_multiplicator => re_multiplicator(438), ---  -0.932983398438
            im_multiplicator => im_multiplicator(438), --- j0.359924316406
            data_re_out => mul_re_out(438),
            data_im_out => mul_im_out(438)
        );

 
    UMUL_439 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(439),
            data_im_in => first_stage_im_out(439),
            re_multiplicator => re_multiplicator(439), ---  -0.863952636719
            im_multiplicator => im_multiplicator(439), --- j0.503540039062
            data_re_out => mul_re_out(439),
            data_im_out => mul_im_out(439)
        );

 
    UMUL_440 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(440),
            data_im_in => first_stage_im_out(440),
            re_multiplicator => re_multiplicator(440), ---  -0.773010253906
            im_multiplicator => im_multiplicator(440), --- j0.634399414062
            data_re_out => mul_re_out(440),
            data_im_out => mul_im_out(440)
        );

 
    UMUL_441 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(441),
            data_im_in => first_stage_im_out(441),
            re_multiplicator => re_multiplicator(441), ---  -0.662414550781
            im_multiplicator => im_multiplicator(441), --- j0.749145507812
            data_re_out => mul_re_out(441),
            data_im_out => mul_im_out(441)
        );

 
    UMUL_442 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(442),
            data_im_in => first_stage_im_out(442),
            re_multiplicator => re_multiplicator(442), ---  -0.534973144531
            im_multiplicator => im_multiplicator(442), --- j0.844848632812
            data_re_out => mul_re_out(442),
            data_im_out => mul_im_out(442)
        );

 
    UMUL_443 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(443),
            data_im_in => first_stage_im_out(443),
            re_multiplicator => re_multiplicator(443), ---  -0.393981933594
            im_multiplicator => im_multiplicator(443), --- j0.919128417969
            data_re_out => mul_re_out(443),
            data_im_out => mul_im_out(443)
        );

 
    UMUL_444 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(444),
            data_im_in => first_stage_im_out(444),
            re_multiplicator => re_multiplicator(444), ---  -0.242980957031
            im_multiplicator => im_multiplicator(444), --- j0.970031738281
            data_re_out => mul_re_out(444),
            data_im_out => mul_im_out(444)
        );

 
    UMUL_445 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(445),
            data_im_in => first_stage_im_out(445),
            re_multiplicator => re_multiplicator(445), ---  -0.0858154296875
            im_multiplicator => im_multiplicator(445), --- j0.996337890625
            data_re_out => mul_re_out(445),
            data_im_out => mul_im_out(445)
        );

 
    UMUL_446 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(446),
            data_im_in => first_stage_im_out(446),
            re_multiplicator => re_multiplicator(446), ---  0.0735473632812
            im_multiplicator => im_multiplicator(446), --- j0.997314453125
            data_re_out => mul_re_out(446),
            data_im_out => mul_im_out(446)
        );

 
    UMUL_447 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(447),
            data_im_in => first_stage_im_out(447),
            re_multiplicator => re_multiplicator(447), ---  0.231079101562
            im_multiplicator => im_multiplicator(447), --- j0.972961425781
            data_re_out => mul_re_out(447),
            data_im_out => mul_im_out(447)
        );

 
    UMUL_448 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(448),
            data_im_in => first_stage_im_out(448),
            data_re_out => mul_re_out(448),
            data_im_out => mul_im_out(448)
        );

 
    UMUL_449 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(449),
            data_im_in => first_stage_im_out(449),
            re_multiplicator => re_multiplicator(449), ---  0.985290527344
            im_multiplicator => im_multiplicator(449), --- j-0.170959472656
            data_re_out => mul_re_out(449),
            data_im_out => mul_im_out(449)
        );

 
    UMUL_450 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(450),
            data_im_in => first_stage_im_out(450),
            re_multiplicator => re_multiplicator(450), ---  0.941528320312
            im_multiplicator => im_multiplicator(450), --- j-0.3369140625
            data_re_out => mul_re_out(450),
            data_im_out => mul_im_out(450)
        );

 
    UMUL_451 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(451),
            data_im_in => first_stage_im_out(451),
            re_multiplicator => re_multiplicator(451), ---  0.8701171875
            im_multiplicator => im_multiplicator(451), --- j-0.492919921875
            data_re_out => mul_re_out(451),
            data_im_out => mul_im_out(451)
        );

 
    UMUL_452 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(452),
            data_im_in => first_stage_im_out(452),
            re_multiplicator => re_multiplicator(452), ---  0.773010253906
            im_multiplicator => im_multiplicator(452), --- j-0.634399414062
            data_re_out => mul_re_out(452),
            data_im_out => mul_im_out(452)
        );

 
    UMUL_453 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(453),
            data_im_in => first_stage_im_out(453),
            re_multiplicator => re_multiplicator(453), ---  0.653198242188
            im_multiplicator => im_multiplicator(453), --- j-0.757202148438
            data_re_out => mul_re_out(453),
            data_im_out => mul_im_out(453)
        );

 
    UMUL_454 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(454),
            data_im_in => first_stage_im_out(454),
            re_multiplicator => re_multiplicator(454), ---  0.514099121094
            im_multiplicator => im_multiplicator(454), --- j-0.857727050781
            data_re_out => mul_re_out(454),
            data_im_out => mul_im_out(454)
        );

 
    UMUL_455 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(455),
            data_im_in => first_stage_im_out(455),
            re_multiplicator => re_multiplicator(455), ---  0.359924316406
            im_multiplicator => im_multiplicator(455), --- j-0.932983398438
            data_re_out => mul_re_out(455),
            data_im_out => mul_im_out(455)
        );

 
    UMUL_456 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(456),
            data_im_in => first_stage_im_out(456),
            re_multiplicator => re_multiplicator(456), ---  0.195068359375
            im_multiplicator => im_multiplicator(456), --- j-0.980773925781
            data_re_out => mul_re_out(456),
            data_im_out => mul_im_out(456)
        );

 
    UMUL_457 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(457),
            data_im_in => first_stage_im_out(457),
            re_multiplicator => re_multiplicator(457), ---  0.0245361328125
            im_multiplicator => im_multiplicator(457), --- j-0.999694824219
            data_re_out => mul_re_out(457),
            data_im_out => mul_im_out(457)
        );

 
    UMUL_458 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(458),
            data_im_in => first_stage_im_out(458),
            re_multiplicator => re_multiplicator(458), ---  -0.146728515625
            im_multiplicator => im_multiplicator(458), --- j-0.989196777344
            data_re_out => mul_re_out(458),
            data_im_out => mul_im_out(458)
        );

 
    UMUL_459 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(459),
            data_im_in => first_stage_im_out(459),
            re_multiplicator => re_multiplicator(459), ---  -0.313659667969
            im_multiplicator => im_multiplicator(459), --- j-0.949523925781
            data_re_out => mul_re_out(459),
            data_im_out => mul_im_out(459)
        );

 
    UMUL_460 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(460),
            data_im_in => first_stage_im_out(460),
            re_multiplicator => re_multiplicator(460), ---  -0.471374511719
            im_multiplicator => im_multiplicator(460), --- j-0.881896972656
            data_re_out => mul_re_out(460),
            data_im_out => mul_im_out(460)
        );

 
    UMUL_461 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(461),
            data_im_in => first_stage_im_out(461),
            re_multiplicator => re_multiplicator(461), ---  -0.615234375
            im_multiplicator => im_multiplicator(461), --- j-0.788330078125
            data_re_out => mul_re_out(461),
            data_im_out => mul_im_out(461)
        );

 
    UMUL_462 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(462),
            data_im_in => first_stage_im_out(462),
            re_multiplicator => re_multiplicator(462), ---  -0.740966796875
            im_multiplicator => im_multiplicator(462), --- j-0.671569824219
            data_re_out => mul_re_out(462),
            data_im_out => mul_im_out(462)
        );

 
    UMUL_463 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(463),
            data_im_in => first_stage_im_out(463),
            re_multiplicator => re_multiplicator(463), ---  -0.844848632812
            im_multiplicator => im_multiplicator(463), --- j-0.534973144531
            data_re_out => mul_re_out(463),
            data_im_out => mul_im_out(463)
        );

 
    UMUL_464 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(464),
            data_im_in => first_stage_im_out(464),
            re_multiplicator => re_multiplicator(464), ---  -0.923889160156
            im_multiplicator => im_multiplicator(464), --- j-0.382690429688
            data_re_out => mul_re_out(464),
            data_im_out => mul_im_out(464)
        );

 
    UMUL_465 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(465),
            data_im_in => first_stage_im_out(465),
            re_multiplicator => re_multiplicator(465), ---  -0.975708007812
            im_multiplicator => im_multiplicator(465), --- j-0.219116210938
            data_re_out => mul_re_out(465),
            data_im_out => mul_im_out(465)
        );

 
    UMUL_466 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(466),
            data_im_in => first_stage_im_out(466),
            re_multiplicator => re_multiplicator(466), ---  -0.998779296875
            im_multiplicator => im_multiplicator(466), --- j-0.049072265625
            data_re_out => mul_re_out(466),
            data_im_out => mul_im_out(466)
        );

 
    UMUL_467 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(467),
            data_im_in => first_stage_im_out(467),
            re_multiplicator => re_multiplicator(467), ---  -0.992492675781
            im_multiplicator => im_multiplicator(467), --- j0.122436523438
            data_re_out => mul_re_out(467),
            data_im_out => mul_im_out(467)
        );

 
    UMUL_468 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(468),
            data_im_in => first_stage_im_out(468),
            re_multiplicator => re_multiplicator(468), ---  -0.956970214844
            im_multiplicator => im_multiplicator(468), --- j0.290283203125
            data_re_out => mul_re_out(468),
            data_im_out => mul_im_out(468)
        );

 
    UMUL_469 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(469),
            data_im_in => first_stage_im_out(469),
            re_multiplicator => re_multiplicator(469), ---  -0.893249511719
            im_multiplicator => im_multiplicator(469), --- j0.449584960938
            data_re_out => mul_re_out(469),
            data_im_out => mul_im_out(469)
        );

 
    UMUL_470 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(470),
            data_im_in => first_stage_im_out(470),
            re_multiplicator => re_multiplicator(470), ---  -0.80322265625
            im_multiplicator => im_multiplicator(470), --- j0.595703125
            data_re_out => mul_re_out(470),
            data_im_out => mul_im_out(470)
        );

 
    UMUL_471 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(471),
            data_im_in => first_stage_im_out(471),
            re_multiplicator => re_multiplicator(471), ---  -0.689514160156
            im_multiplicator => im_multiplicator(471), --- j0.724243164062
            data_re_out => mul_re_out(471),
            data_im_out => mul_im_out(471)
        );

 
    UMUL_472 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(472),
            data_im_in => first_stage_im_out(472),
            re_multiplicator => re_multiplicator(472), ---  -0.555541992188
            im_multiplicator => im_multiplicator(472), --- j0.831481933594
            data_re_out => mul_re_out(472),
            data_im_out => mul_im_out(472)
        );

 
    UMUL_473 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(473),
            data_im_in => first_stage_im_out(473),
            re_multiplicator => re_multiplicator(473), ---  -0.405212402344
            im_multiplicator => im_multiplicator(473), --- j0.914184570312
            data_re_out => mul_re_out(473),
            data_im_out => mul_im_out(473)
        );

 
    UMUL_474 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(474),
            data_im_in => first_stage_im_out(474),
            re_multiplicator => re_multiplicator(474), ---  -0.242980957031
            im_multiplicator => im_multiplicator(474), --- j0.970031738281
            data_re_out => mul_re_out(474),
            data_im_out => mul_im_out(474)
        );

 
    UMUL_475 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(475),
            data_im_in => first_stage_im_out(475),
            re_multiplicator => re_multiplicator(475), ---  -0.0735473632812
            im_multiplicator => im_multiplicator(475), --- j0.997314453125
            data_re_out => mul_re_out(475),
            data_im_out => mul_im_out(475)
        );

 
    UMUL_476 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(476),
            data_im_in => first_stage_im_out(476),
            re_multiplicator => re_multiplicator(476), ---  0.0980224609375
            im_multiplicator => im_multiplicator(476), --- j0.995178222656
            data_re_out => mul_re_out(476),
            data_im_out => mul_im_out(476)
        );

 
    UMUL_477 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(477),
            data_im_in => first_stage_im_out(477),
            re_multiplicator => re_multiplicator(477), ---  0.266723632812
            im_multiplicator => im_multiplicator(477), --- j0.963806152344
            data_re_out => mul_re_out(477),
            data_im_out => mul_im_out(477)
        );

 
    UMUL_478 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(478),
            data_im_in => first_stage_im_out(478),
            re_multiplicator => re_multiplicator(478), ---  0.427551269531
            im_multiplicator => im_multiplicator(478), --- j0.903991699219
            data_re_out => mul_re_out(478),
            data_im_out => mul_im_out(478)
        );

 
    UMUL_479 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(479),
            data_im_in => first_stage_im_out(479),
            re_multiplicator => re_multiplicator(479), ---  0.575805664062
            im_multiplicator => im_multiplicator(479), --- j0.817565917969
            data_re_out => mul_re_out(479),
            data_im_out => mul_im_out(479)
        );

 
    UMUL_480 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(480),
            data_im_in => first_stage_im_out(480),
            data_re_out => mul_re_out(480),
            data_im_out => mul_im_out(480)
        );

 
    UMUL_481 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(481),
            data_im_in => first_stage_im_out(481),
            re_multiplicator => re_multiplicator(481), ---  0.983093261719
            im_multiplicator => im_multiplicator(481), --- j-0.183044433594
            data_re_out => mul_re_out(481),
            data_im_out => mul_im_out(481)
        );

 
    UMUL_482 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(482),
            data_im_in => first_stage_im_out(482),
            re_multiplicator => re_multiplicator(482), ---  0.932983398438
            im_multiplicator => im_multiplicator(482), --- j-0.359924316406
            data_re_out => mul_re_out(482),
            data_im_out => mul_im_out(482)
        );

 
    UMUL_483 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(483),
            data_im_in => first_stage_im_out(483),
            re_multiplicator => re_multiplicator(483), ---  0.851379394531
            im_multiplicator => im_multiplicator(483), --- j-0.524597167969
            data_re_out => mul_re_out(483),
            data_im_out => mul_im_out(483)
        );

 
    UMUL_484 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(484),
            data_im_in => first_stage_im_out(484),
            re_multiplicator => re_multiplicator(484), ---  0.740966796875
            im_multiplicator => im_multiplicator(484), --- j-0.671569824219
            data_re_out => mul_re_out(484),
            data_im_out => mul_im_out(484)
        );

 
    UMUL_485 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(485),
            data_im_in => first_stage_im_out(485),
            re_multiplicator => re_multiplicator(485), ---  0.605529785156
            im_multiplicator => im_multiplicator(485), --- j-0.795837402344
            data_re_out => mul_re_out(485),
            data_im_out => mul_im_out(485)
        );

 
    UMUL_486 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(486),
            data_im_in => first_stage_im_out(486),
            re_multiplicator => re_multiplicator(486), ---  0.449584960938
            im_multiplicator => im_multiplicator(486), --- j-0.893249511719
            data_re_out => mul_re_out(486),
            data_im_out => mul_im_out(486)
        );

 
    UMUL_487 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(487),
            data_im_in => first_stage_im_out(487),
            re_multiplicator => re_multiplicator(487), ---  0.278503417969
            im_multiplicator => im_multiplicator(487), --- j-0.96044921875
            data_re_out => mul_re_out(487),
            data_im_out => mul_im_out(487)
        );

 
    UMUL_488 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(488),
            data_im_in => first_stage_im_out(488),
            re_multiplicator => re_multiplicator(488), ---  0.0980224609375
            im_multiplicator => im_multiplicator(488), --- j-0.995178222656
            data_re_out => mul_re_out(488),
            data_im_out => mul_im_out(488)
        );

 
    UMUL_489 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(489),
            data_im_in => first_stage_im_out(489),
            re_multiplicator => re_multiplicator(489), ---  -0.0858154296875
            im_multiplicator => im_multiplicator(489), --- j-0.996337890625
            data_re_out => mul_re_out(489),
            data_im_out => mul_im_out(489)
        );

 
    UMUL_490 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(490),
            data_im_in => first_stage_im_out(490),
            re_multiplicator => re_multiplicator(490), ---  -0.266723632812
            im_multiplicator => im_multiplicator(490), --- j-0.963806152344
            data_re_out => mul_re_out(490),
            data_im_out => mul_im_out(490)
        );

 
    UMUL_491 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(491),
            data_im_in => first_stage_im_out(491),
            re_multiplicator => re_multiplicator(491), ---  -0.438598632812
            im_multiplicator => im_multiplicator(491), --- j-0.898681640625
            data_re_out => mul_re_out(491),
            data_im_out => mul_im_out(491)
        );

 
    UMUL_492 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(492),
            data_im_in => first_stage_im_out(492),
            re_multiplicator => re_multiplicator(492), ---  -0.595703125
            im_multiplicator => im_multiplicator(492), --- j-0.80322265625
            data_re_out => mul_re_out(492),
            data_im_out => mul_im_out(492)
        );

 
    UMUL_493 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(493),
            data_im_in => first_stage_im_out(493),
            re_multiplicator => re_multiplicator(493), ---  -0.732666015625
            im_multiplicator => im_multiplicator(493), --- j-0.680603027344
            data_re_out => mul_re_out(493),
            data_im_out => mul_im_out(493)
        );

 
    UMUL_494 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(494),
            data_im_in => first_stage_im_out(494),
            re_multiplicator => re_multiplicator(494), ---  -0.844848632812
            im_multiplicator => im_multiplicator(494), --- j-0.534973144531
            data_re_out => mul_re_out(494),
            data_im_out => mul_im_out(494)
        );

 
    UMUL_495 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(495),
            data_im_in => first_stage_im_out(495),
            re_multiplicator => re_multiplicator(495), ---  -0.928527832031
            im_multiplicator => im_multiplicator(495), --- j-0.371337890625
            data_re_out => mul_re_out(495),
            data_im_out => mul_im_out(495)
        );

 
    UMUL_496 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(496),
            data_im_in => first_stage_im_out(496),
            re_multiplicator => re_multiplicator(496), ---  -0.980773925781
            im_multiplicator => im_multiplicator(496), --- j-0.195068359375
            data_re_out => mul_re_out(496),
            data_im_out => mul_im_out(496)
        );

 
    UMUL_497 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(497),
            data_im_in => first_stage_im_out(497),
            re_multiplicator => re_multiplicator(497), ---  -0.999938964844
            im_multiplicator => im_multiplicator(497), --- j-0.0122680664062
            data_re_out => mul_re_out(497),
            data_im_out => mul_im_out(497)
        );

 
    UMUL_498 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(498),
            data_im_in => first_stage_im_out(498),
            re_multiplicator => re_multiplicator(498), ---  -0.985290527344
            im_multiplicator => im_multiplicator(498), --- j0.170959472656
            data_re_out => mul_re_out(498),
            data_im_out => mul_im_out(498)
        );

 
    UMUL_499 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(499),
            data_im_in => first_stage_im_out(499),
            re_multiplicator => re_multiplicator(499), ---  -0.937316894531
            im_multiplicator => im_multiplicator(499), --- j0.348388671875
            data_re_out => mul_re_out(499),
            data_im_out => mul_im_out(499)
        );

 
    UMUL_500 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(500),
            data_im_in => first_stage_im_out(500),
            re_multiplicator => re_multiplicator(500), ---  -0.857727050781
            im_multiplicator => im_multiplicator(500), --- j0.514099121094
            data_re_out => mul_re_out(500),
            data_im_out => mul_im_out(500)
        );

 
    UMUL_501 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(501),
            data_im_in => first_stage_im_out(501),
            re_multiplicator => re_multiplicator(501), ---  -0.749145507812
            im_multiplicator => im_multiplicator(501), --- j0.662414550781
            data_re_out => mul_re_out(501),
            data_im_out => mul_im_out(501)
        );

 
    UMUL_502 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(502),
            data_im_in => first_stage_im_out(502),
            re_multiplicator => re_multiplicator(502), ---  -0.615234375
            im_multiplicator => im_multiplicator(502), --- j0.788330078125
            data_re_out => mul_re_out(502),
            data_im_out => mul_im_out(502)
        );

 
    UMUL_503 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(503),
            data_im_in => first_stage_im_out(503),
            re_multiplicator => re_multiplicator(503), ---  -0.460510253906
            im_multiplicator => im_multiplicator(503), --- j0.887634277344
            data_re_out => mul_re_out(503),
            data_im_out => mul_im_out(503)
        );

 
    UMUL_504 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(504),
            data_im_in => first_stage_im_out(504),
            re_multiplicator => re_multiplicator(504), ---  -0.290283203125
            im_multiplicator => im_multiplicator(504), --- j0.956970214844
            data_re_out => mul_re_out(504),
            data_im_out => mul_im_out(504)
        );

 
    UMUL_505 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(505),
            data_im_in => first_stage_im_out(505),
            re_multiplicator => re_multiplicator(505), ---  -0.110229492188
            im_multiplicator => im_multiplicator(505), --- j0.993896484375
            data_re_out => mul_re_out(505),
            data_im_out => mul_im_out(505)
        );

 
    UMUL_506 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(506),
            data_im_in => first_stage_im_out(506),
            re_multiplicator => re_multiplicator(506), ---  0.0735473632812
            im_multiplicator => im_multiplicator(506), --- j0.997314453125
            data_re_out => mul_re_out(506),
            data_im_out => mul_im_out(506)
        );

 
    UMUL_507 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(507),
            data_im_in => first_stage_im_out(507),
            re_multiplicator => re_multiplicator(507), ---  0.2548828125
            im_multiplicator => im_multiplicator(507), --- j0.966979980469
            data_re_out => mul_re_out(507),
            data_im_out => mul_im_out(507)
        );

 
    UMUL_508 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(508),
            data_im_in => first_stage_im_out(508),
            re_multiplicator => re_multiplicator(508), ---  0.427551269531
            im_multiplicator => im_multiplicator(508), --- j0.903991699219
            data_re_out => mul_re_out(508),
            data_im_out => mul_im_out(508)
        );

 
    UMUL_509 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(509),
            data_im_in => first_stage_im_out(509),
            re_multiplicator => re_multiplicator(509), ---  0.585815429688
            im_multiplicator => im_multiplicator(509), --- j0.810485839844
            data_re_out => mul_re_out(509),
            data_im_out => mul_im_out(509)
        );

 
    UMUL_510 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(510),
            data_im_in => first_stage_im_out(510),
            re_multiplicator => re_multiplicator(510), ---  0.724243164062
            im_multiplicator => im_multiplicator(510), --- j0.689514160156
            data_re_out => mul_re_out(510),
            data_im_out => mul_im_out(510)
        );

 
    UMUL_511 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(511),
            data_im_in => first_stage_im_out(511),
            re_multiplicator => re_multiplicator(511), ---  0.838195800781
            im_multiplicator => im_multiplicator(511), --- j0.545349121094
            data_re_out => mul_re_out(511),
            data_im_out => mul_im_out(511)
        );

end Behavioral;
