library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity fft_pt512 is
    GENERIC (
        ctrl_start     : INTEGER := 0
    );
    PORT (
        tmp_first_stage_re_out, tmp_first_stage_im_out: OUT STD_LOGIC_VECTOR(511 DOWNTO 0);
        tmp_mul_re_out, tmp_mul_im_out : OUT STD_LOGIC_VECTOR(511 DOWNTO 0);

        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        bypass         : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
        ctrl_delay     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

        data_re_in     : IN STD_LOGIC_VECTOR(511 DOWNTO 0);
        data_im_in     : IN STD_LOGIC_VECTOR(511 DOWNTO 0);

        data_re_out    : OUT STD_LOGIC_VECTOR(511 DOWNTO 0);
        data_im_out    : OUT STD_LOGIC_VECTOR(511 DOWNTO 0)
    );
end fft_pt512;

architecture Behavioral of fft_pt512 is

component fft_pt16 is
    GENERIC (
        ctrl_start     : INTEGER
    );
    PORT (
        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        bypass         : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        ctrl_delay     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

        data_re_in     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_im_in     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

        data_re_out    : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_im_out    : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
end component;

component fft_pt32 is
    GENERIC (
        ctrl_start       : INTEGER
    );
    PORT (
        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        bypass         : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        ctrl_delay     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);

        data_re_in     : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        data_im_in     : IN STD_LOGIC_VECTOR(31 DOWNTO 0);

        data_re_out     : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        data_im_out     : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
end component;

component complex_multiplier is
    GENERIC (
        ctrl_start       : INTEGER
    );
    PORT (
        clk              : IN STD_LOGIC;
        rst              : IN STD_LOGIC;
        ce               : IN STD_LOGIC;
        bypass           : IN STD_LOGIC;
        ctrl_delay       : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_in       : IN STD_LOGIC;
        data_im_in       : IN STD_LOGIC;
        re_multiplicator : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        im_multiplicator : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_out      : OUT STD_LOGIC;
        data_im_out      : OUT STD_LOGIC
    );
end component;

component multiplier_mul1 IS
    GENERIC (
        ctrl_start : INTEGER := 0
    );
    PORT (
        clk             : IN STD_LOGIC;
        rst             : IN STD_LOGIC;
        ce              : IN STD_LOGIC;
        bypass          : IN STD_LOGIC;
        ctrl_delay      : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_in      : IN STD_LOGIC;
        data_im_in      : IN STD_LOGIC;
        data_re_out     : OUT STD_LOGIC;
        data_im_out     : OUT STD_LOGIC
    );
END component;

component multiplier_mulminusj IS
    GENERIC (
        ctrl_start : INTEGER := 0
    );
    PORT (
        clk             : IN STD_LOGIC;
        rst             : IN STD_LOGIC;
        ce              : IN STD_LOGIC;
        bypass          : IN STD_LOGIC;
        ctrl_delay      : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        data_re_in      : IN STD_LOGIC;
        data_im_in      : IN STD_LOGIC;
        data_re_out     : OUT STD_LOGIC;
        data_im_out     : OUT STD_LOGIC
    );
END component;

COMPONENT Dff_regN_Nout IS
    GENERIC (N : INTEGER);
    PORT (  
        D      : IN STD_LOGIC;
        clk    : IN STD_LOGIC;
        Q      : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        QN     : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0)
    );
END COMPONENT;

signal first_stage_re_out, first_stage_im_out: STD_LOGIC_VECTOR(511 DOWNTO 0);
signal mul_re_out, mul_im_out : STD_LOGIC_VECTOR(511 DOWNTO 0);


begin

    tmp_first_stage_re_out <= first_stage_re_out;
    tmp_first_stage_im_out <= first_stage_im_out;
    tmp_mul_re_out <= mul_re_out;
    tmp_mul_im_out <= mul_im_out;

    --- left-hand-side processors
    ULFFT_PT16_0 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(0),
            data_re_in(1) => data_re_in(32),
            data_re_in(2) => data_re_in(64),
            data_re_in(3) => data_re_in(96),
            data_re_in(4) => data_re_in(128),
            data_re_in(5) => data_re_in(160),
            data_re_in(6) => data_re_in(192),
            data_re_in(7) => data_re_in(224),
            data_re_in(8) => data_re_in(256),
            data_re_in(9) => data_re_in(288),
            data_re_in(10) => data_re_in(320),
            data_re_in(11) => data_re_in(352),
            data_re_in(12) => data_re_in(384),
            data_re_in(13) => data_re_in(416),
            data_re_in(14) => data_re_in(448),
            data_re_in(15) => data_re_in(480),
            data_im_in(0) => data_im_in(0),
            data_im_in(1) => data_im_in(32),
            data_im_in(2) => data_im_in(64),
            data_im_in(3) => data_im_in(96),
            data_im_in(4) => data_im_in(128),
            data_im_in(5) => data_im_in(160),
            data_im_in(6) => data_im_in(192),
            data_im_in(7) => data_im_in(224),
            data_im_in(8) => data_im_in(256),
            data_im_in(9) => data_im_in(288),
            data_im_in(10) => data_im_in(320),
            data_im_in(11) => data_im_in(352),
            data_im_in(12) => data_im_in(384),
            data_im_in(13) => data_im_in(416),
            data_im_in(14) => data_im_in(448),
            data_im_in(15) => data_im_in(480),
            data_re_out(0) => first_stage_re_out(0),
            data_re_out(1) => first_stage_re_out(32),
            data_re_out(2) => first_stage_re_out(64),
            data_re_out(3) => first_stage_re_out(96),
            data_re_out(4) => first_stage_re_out(128),
            data_re_out(5) => first_stage_re_out(160),
            data_re_out(6) => first_stage_re_out(192),
            data_re_out(7) => first_stage_re_out(224),
            data_re_out(8) => first_stage_re_out(256),
            data_re_out(9) => first_stage_re_out(288),
            data_re_out(10) => first_stage_re_out(320),
            data_re_out(11) => first_stage_re_out(352),
            data_re_out(12) => first_stage_re_out(384),
            data_re_out(13) => first_stage_re_out(416),
            data_re_out(14) => first_stage_re_out(448),
            data_re_out(15) => first_stage_re_out(480),
            data_im_out(0) => first_stage_im_out(0),
            data_im_out(1) => first_stage_im_out(32),
            data_im_out(2) => first_stage_im_out(64),
            data_im_out(3) => first_stage_im_out(96),
            data_im_out(4) => first_stage_im_out(128),
            data_im_out(5) => first_stage_im_out(160),
            data_im_out(6) => first_stage_im_out(192),
            data_im_out(7) => first_stage_im_out(224),
            data_im_out(8) => first_stage_im_out(256),
            data_im_out(9) => first_stage_im_out(288),
            data_im_out(10) => first_stage_im_out(320),
            data_im_out(11) => first_stage_im_out(352),
            data_im_out(12) => first_stage_im_out(384),
            data_im_out(13) => first_stage_im_out(416),
            data_im_out(14) => first_stage_im_out(448),
            data_im_out(15) => first_stage_im_out(480)
        );

    ULFFT_PT16_1 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(1),
            data_re_in(1) => data_re_in(33),
            data_re_in(2) => data_re_in(65),
            data_re_in(3) => data_re_in(97),
            data_re_in(4) => data_re_in(129),
            data_re_in(5) => data_re_in(161),
            data_re_in(6) => data_re_in(193),
            data_re_in(7) => data_re_in(225),
            data_re_in(8) => data_re_in(257),
            data_re_in(9) => data_re_in(289),
            data_re_in(10) => data_re_in(321),
            data_re_in(11) => data_re_in(353),
            data_re_in(12) => data_re_in(385),
            data_re_in(13) => data_re_in(417),
            data_re_in(14) => data_re_in(449),
            data_re_in(15) => data_re_in(481),
            data_im_in(0) => data_im_in(1),
            data_im_in(1) => data_im_in(33),
            data_im_in(2) => data_im_in(65),
            data_im_in(3) => data_im_in(97),
            data_im_in(4) => data_im_in(129),
            data_im_in(5) => data_im_in(161),
            data_im_in(6) => data_im_in(193),
            data_im_in(7) => data_im_in(225),
            data_im_in(8) => data_im_in(257),
            data_im_in(9) => data_im_in(289),
            data_im_in(10) => data_im_in(321),
            data_im_in(11) => data_im_in(353),
            data_im_in(12) => data_im_in(385),
            data_im_in(13) => data_im_in(417),
            data_im_in(14) => data_im_in(449),
            data_im_in(15) => data_im_in(481),
            data_re_out(0) => first_stage_re_out(1),
            data_re_out(1) => first_stage_re_out(33),
            data_re_out(2) => first_stage_re_out(65),
            data_re_out(3) => first_stage_re_out(97),
            data_re_out(4) => first_stage_re_out(129),
            data_re_out(5) => first_stage_re_out(161),
            data_re_out(6) => first_stage_re_out(193),
            data_re_out(7) => first_stage_re_out(225),
            data_re_out(8) => first_stage_re_out(257),
            data_re_out(9) => first_stage_re_out(289),
            data_re_out(10) => first_stage_re_out(321),
            data_re_out(11) => first_stage_re_out(353),
            data_re_out(12) => first_stage_re_out(385),
            data_re_out(13) => first_stage_re_out(417),
            data_re_out(14) => first_stage_re_out(449),
            data_re_out(15) => first_stage_re_out(481),
            data_im_out(0) => first_stage_im_out(1),
            data_im_out(1) => first_stage_im_out(33),
            data_im_out(2) => first_stage_im_out(65),
            data_im_out(3) => first_stage_im_out(97),
            data_im_out(4) => first_stage_im_out(129),
            data_im_out(5) => first_stage_im_out(161),
            data_im_out(6) => first_stage_im_out(193),
            data_im_out(7) => first_stage_im_out(225),
            data_im_out(8) => first_stage_im_out(257),
            data_im_out(9) => first_stage_im_out(289),
            data_im_out(10) => first_stage_im_out(321),
            data_im_out(11) => first_stage_im_out(353),
            data_im_out(12) => first_stage_im_out(385),
            data_im_out(13) => first_stage_im_out(417),
            data_im_out(14) => first_stage_im_out(449),
            data_im_out(15) => first_stage_im_out(481)
        );

    ULFFT_PT16_2 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(2),
            data_re_in(1) => data_re_in(34),
            data_re_in(2) => data_re_in(66),
            data_re_in(3) => data_re_in(98),
            data_re_in(4) => data_re_in(130),
            data_re_in(5) => data_re_in(162),
            data_re_in(6) => data_re_in(194),
            data_re_in(7) => data_re_in(226),
            data_re_in(8) => data_re_in(258),
            data_re_in(9) => data_re_in(290),
            data_re_in(10) => data_re_in(322),
            data_re_in(11) => data_re_in(354),
            data_re_in(12) => data_re_in(386),
            data_re_in(13) => data_re_in(418),
            data_re_in(14) => data_re_in(450),
            data_re_in(15) => data_re_in(482),
            data_im_in(0) => data_im_in(2),
            data_im_in(1) => data_im_in(34),
            data_im_in(2) => data_im_in(66),
            data_im_in(3) => data_im_in(98),
            data_im_in(4) => data_im_in(130),
            data_im_in(5) => data_im_in(162),
            data_im_in(6) => data_im_in(194),
            data_im_in(7) => data_im_in(226),
            data_im_in(8) => data_im_in(258),
            data_im_in(9) => data_im_in(290),
            data_im_in(10) => data_im_in(322),
            data_im_in(11) => data_im_in(354),
            data_im_in(12) => data_im_in(386),
            data_im_in(13) => data_im_in(418),
            data_im_in(14) => data_im_in(450),
            data_im_in(15) => data_im_in(482),
            data_re_out(0) => first_stage_re_out(2),
            data_re_out(1) => first_stage_re_out(34),
            data_re_out(2) => first_stage_re_out(66),
            data_re_out(3) => first_stage_re_out(98),
            data_re_out(4) => first_stage_re_out(130),
            data_re_out(5) => first_stage_re_out(162),
            data_re_out(6) => first_stage_re_out(194),
            data_re_out(7) => first_stage_re_out(226),
            data_re_out(8) => first_stage_re_out(258),
            data_re_out(9) => first_stage_re_out(290),
            data_re_out(10) => first_stage_re_out(322),
            data_re_out(11) => first_stage_re_out(354),
            data_re_out(12) => first_stage_re_out(386),
            data_re_out(13) => first_stage_re_out(418),
            data_re_out(14) => first_stage_re_out(450),
            data_re_out(15) => first_stage_re_out(482),
            data_im_out(0) => first_stage_im_out(2),
            data_im_out(1) => first_stage_im_out(34),
            data_im_out(2) => first_stage_im_out(66),
            data_im_out(3) => first_stage_im_out(98),
            data_im_out(4) => first_stage_im_out(130),
            data_im_out(5) => first_stage_im_out(162),
            data_im_out(6) => first_stage_im_out(194),
            data_im_out(7) => first_stage_im_out(226),
            data_im_out(8) => first_stage_im_out(258),
            data_im_out(9) => first_stage_im_out(290),
            data_im_out(10) => first_stage_im_out(322),
            data_im_out(11) => first_stage_im_out(354),
            data_im_out(12) => first_stage_im_out(386),
            data_im_out(13) => first_stage_im_out(418),
            data_im_out(14) => first_stage_im_out(450),
            data_im_out(15) => first_stage_im_out(482)
        );

    ULFFT_PT16_3 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(3),
            data_re_in(1) => data_re_in(35),
            data_re_in(2) => data_re_in(67),
            data_re_in(3) => data_re_in(99),
            data_re_in(4) => data_re_in(131),
            data_re_in(5) => data_re_in(163),
            data_re_in(6) => data_re_in(195),
            data_re_in(7) => data_re_in(227),
            data_re_in(8) => data_re_in(259),
            data_re_in(9) => data_re_in(291),
            data_re_in(10) => data_re_in(323),
            data_re_in(11) => data_re_in(355),
            data_re_in(12) => data_re_in(387),
            data_re_in(13) => data_re_in(419),
            data_re_in(14) => data_re_in(451),
            data_re_in(15) => data_re_in(483),
            data_im_in(0) => data_im_in(3),
            data_im_in(1) => data_im_in(35),
            data_im_in(2) => data_im_in(67),
            data_im_in(3) => data_im_in(99),
            data_im_in(4) => data_im_in(131),
            data_im_in(5) => data_im_in(163),
            data_im_in(6) => data_im_in(195),
            data_im_in(7) => data_im_in(227),
            data_im_in(8) => data_im_in(259),
            data_im_in(9) => data_im_in(291),
            data_im_in(10) => data_im_in(323),
            data_im_in(11) => data_im_in(355),
            data_im_in(12) => data_im_in(387),
            data_im_in(13) => data_im_in(419),
            data_im_in(14) => data_im_in(451),
            data_im_in(15) => data_im_in(483),
            data_re_out(0) => first_stage_re_out(3),
            data_re_out(1) => first_stage_re_out(35),
            data_re_out(2) => first_stage_re_out(67),
            data_re_out(3) => first_stage_re_out(99),
            data_re_out(4) => first_stage_re_out(131),
            data_re_out(5) => first_stage_re_out(163),
            data_re_out(6) => first_stage_re_out(195),
            data_re_out(7) => first_stage_re_out(227),
            data_re_out(8) => first_stage_re_out(259),
            data_re_out(9) => first_stage_re_out(291),
            data_re_out(10) => first_stage_re_out(323),
            data_re_out(11) => first_stage_re_out(355),
            data_re_out(12) => first_stage_re_out(387),
            data_re_out(13) => first_stage_re_out(419),
            data_re_out(14) => first_stage_re_out(451),
            data_re_out(15) => first_stage_re_out(483),
            data_im_out(0) => first_stage_im_out(3),
            data_im_out(1) => first_stage_im_out(35),
            data_im_out(2) => first_stage_im_out(67),
            data_im_out(3) => first_stage_im_out(99),
            data_im_out(4) => first_stage_im_out(131),
            data_im_out(5) => first_stage_im_out(163),
            data_im_out(6) => first_stage_im_out(195),
            data_im_out(7) => first_stage_im_out(227),
            data_im_out(8) => first_stage_im_out(259),
            data_im_out(9) => first_stage_im_out(291),
            data_im_out(10) => first_stage_im_out(323),
            data_im_out(11) => first_stage_im_out(355),
            data_im_out(12) => first_stage_im_out(387),
            data_im_out(13) => first_stage_im_out(419),
            data_im_out(14) => first_stage_im_out(451),
            data_im_out(15) => first_stage_im_out(483)
        );

    ULFFT_PT16_4 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(4),
            data_re_in(1) => data_re_in(36),
            data_re_in(2) => data_re_in(68),
            data_re_in(3) => data_re_in(100),
            data_re_in(4) => data_re_in(132),
            data_re_in(5) => data_re_in(164),
            data_re_in(6) => data_re_in(196),
            data_re_in(7) => data_re_in(228),
            data_re_in(8) => data_re_in(260),
            data_re_in(9) => data_re_in(292),
            data_re_in(10) => data_re_in(324),
            data_re_in(11) => data_re_in(356),
            data_re_in(12) => data_re_in(388),
            data_re_in(13) => data_re_in(420),
            data_re_in(14) => data_re_in(452),
            data_re_in(15) => data_re_in(484),
            data_im_in(0) => data_im_in(4),
            data_im_in(1) => data_im_in(36),
            data_im_in(2) => data_im_in(68),
            data_im_in(3) => data_im_in(100),
            data_im_in(4) => data_im_in(132),
            data_im_in(5) => data_im_in(164),
            data_im_in(6) => data_im_in(196),
            data_im_in(7) => data_im_in(228),
            data_im_in(8) => data_im_in(260),
            data_im_in(9) => data_im_in(292),
            data_im_in(10) => data_im_in(324),
            data_im_in(11) => data_im_in(356),
            data_im_in(12) => data_im_in(388),
            data_im_in(13) => data_im_in(420),
            data_im_in(14) => data_im_in(452),
            data_im_in(15) => data_im_in(484),
            data_re_out(0) => first_stage_re_out(4),
            data_re_out(1) => first_stage_re_out(36),
            data_re_out(2) => first_stage_re_out(68),
            data_re_out(3) => first_stage_re_out(100),
            data_re_out(4) => first_stage_re_out(132),
            data_re_out(5) => first_stage_re_out(164),
            data_re_out(6) => first_stage_re_out(196),
            data_re_out(7) => first_stage_re_out(228),
            data_re_out(8) => first_stage_re_out(260),
            data_re_out(9) => first_stage_re_out(292),
            data_re_out(10) => first_stage_re_out(324),
            data_re_out(11) => first_stage_re_out(356),
            data_re_out(12) => first_stage_re_out(388),
            data_re_out(13) => first_stage_re_out(420),
            data_re_out(14) => first_stage_re_out(452),
            data_re_out(15) => first_stage_re_out(484),
            data_im_out(0) => first_stage_im_out(4),
            data_im_out(1) => first_stage_im_out(36),
            data_im_out(2) => first_stage_im_out(68),
            data_im_out(3) => first_stage_im_out(100),
            data_im_out(4) => first_stage_im_out(132),
            data_im_out(5) => first_stage_im_out(164),
            data_im_out(6) => first_stage_im_out(196),
            data_im_out(7) => first_stage_im_out(228),
            data_im_out(8) => first_stage_im_out(260),
            data_im_out(9) => first_stage_im_out(292),
            data_im_out(10) => first_stage_im_out(324),
            data_im_out(11) => first_stage_im_out(356),
            data_im_out(12) => first_stage_im_out(388),
            data_im_out(13) => first_stage_im_out(420),
            data_im_out(14) => first_stage_im_out(452),
            data_im_out(15) => first_stage_im_out(484)
        );

    ULFFT_PT16_5 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(5),
            data_re_in(1) => data_re_in(37),
            data_re_in(2) => data_re_in(69),
            data_re_in(3) => data_re_in(101),
            data_re_in(4) => data_re_in(133),
            data_re_in(5) => data_re_in(165),
            data_re_in(6) => data_re_in(197),
            data_re_in(7) => data_re_in(229),
            data_re_in(8) => data_re_in(261),
            data_re_in(9) => data_re_in(293),
            data_re_in(10) => data_re_in(325),
            data_re_in(11) => data_re_in(357),
            data_re_in(12) => data_re_in(389),
            data_re_in(13) => data_re_in(421),
            data_re_in(14) => data_re_in(453),
            data_re_in(15) => data_re_in(485),
            data_im_in(0) => data_im_in(5),
            data_im_in(1) => data_im_in(37),
            data_im_in(2) => data_im_in(69),
            data_im_in(3) => data_im_in(101),
            data_im_in(4) => data_im_in(133),
            data_im_in(5) => data_im_in(165),
            data_im_in(6) => data_im_in(197),
            data_im_in(7) => data_im_in(229),
            data_im_in(8) => data_im_in(261),
            data_im_in(9) => data_im_in(293),
            data_im_in(10) => data_im_in(325),
            data_im_in(11) => data_im_in(357),
            data_im_in(12) => data_im_in(389),
            data_im_in(13) => data_im_in(421),
            data_im_in(14) => data_im_in(453),
            data_im_in(15) => data_im_in(485),
            data_re_out(0) => first_stage_re_out(5),
            data_re_out(1) => first_stage_re_out(37),
            data_re_out(2) => first_stage_re_out(69),
            data_re_out(3) => first_stage_re_out(101),
            data_re_out(4) => first_stage_re_out(133),
            data_re_out(5) => first_stage_re_out(165),
            data_re_out(6) => first_stage_re_out(197),
            data_re_out(7) => first_stage_re_out(229),
            data_re_out(8) => first_stage_re_out(261),
            data_re_out(9) => first_stage_re_out(293),
            data_re_out(10) => first_stage_re_out(325),
            data_re_out(11) => first_stage_re_out(357),
            data_re_out(12) => first_stage_re_out(389),
            data_re_out(13) => first_stage_re_out(421),
            data_re_out(14) => first_stage_re_out(453),
            data_re_out(15) => first_stage_re_out(485),
            data_im_out(0) => first_stage_im_out(5),
            data_im_out(1) => first_stage_im_out(37),
            data_im_out(2) => first_stage_im_out(69),
            data_im_out(3) => first_stage_im_out(101),
            data_im_out(4) => first_stage_im_out(133),
            data_im_out(5) => first_stage_im_out(165),
            data_im_out(6) => first_stage_im_out(197),
            data_im_out(7) => first_stage_im_out(229),
            data_im_out(8) => first_stage_im_out(261),
            data_im_out(9) => first_stage_im_out(293),
            data_im_out(10) => first_stage_im_out(325),
            data_im_out(11) => first_stage_im_out(357),
            data_im_out(12) => first_stage_im_out(389),
            data_im_out(13) => first_stage_im_out(421),
            data_im_out(14) => first_stage_im_out(453),
            data_im_out(15) => first_stage_im_out(485)
        );

    ULFFT_PT16_6 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(6),
            data_re_in(1) => data_re_in(38),
            data_re_in(2) => data_re_in(70),
            data_re_in(3) => data_re_in(102),
            data_re_in(4) => data_re_in(134),
            data_re_in(5) => data_re_in(166),
            data_re_in(6) => data_re_in(198),
            data_re_in(7) => data_re_in(230),
            data_re_in(8) => data_re_in(262),
            data_re_in(9) => data_re_in(294),
            data_re_in(10) => data_re_in(326),
            data_re_in(11) => data_re_in(358),
            data_re_in(12) => data_re_in(390),
            data_re_in(13) => data_re_in(422),
            data_re_in(14) => data_re_in(454),
            data_re_in(15) => data_re_in(486),
            data_im_in(0) => data_im_in(6),
            data_im_in(1) => data_im_in(38),
            data_im_in(2) => data_im_in(70),
            data_im_in(3) => data_im_in(102),
            data_im_in(4) => data_im_in(134),
            data_im_in(5) => data_im_in(166),
            data_im_in(6) => data_im_in(198),
            data_im_in(7) => data_im_in(230),
            data_im_in(8) => data_im_in(262),
            data_im_in(9) => data_im_in(294),
            data_im_in(10) => data_im_in(326),
            data_im_in(11) => data_im_in(358),
            data_im_in(12) => data_im_in(390),
            data_im_in(13) => data_im_in(422),
            data_im_in(14) => data_im_in(454),
            data_im_in(15) => data_im_in(486),
            data_re_out(0) => first_stage_re_out(6),
            data_re_out(1) => first_stage_re_out(38),
            data_re_out(2) => first_stage_re_out(70),
            data_re_out(3) => first_stage_re_out(102),
            data_re_out(4) => first_stage_re_out(134),
            data_re_out(5) => first_stage_re_out(166),
            data_re_out(6) => first_stage_re_out(198),
            data_re_out(7) => first_stage_re_out(230),
            data_re_out(8) => first_stage_re_out(262),
            data_re_out(9) => first_stage_re_out(294),
            data_re_out(10) => first_stage_re_out(326),
            data_re_out(11) => first_stage_re_out(358),
            data_re_out(12) => first_stage_re_out(390),
            data_re_out(13) => first_stage_re_out(422),
            data_re_out(14) => first_stage_re_out(454),
            data_re_out(15) => first_stage_re_out(486),
            data_im_out(0) => first_stage_im_out(6),
            data_im_out(1) => first_stage_im_out(38),
            data_im_out(2) => first_stage_im_out(70),
            data_im_out(3) => first_stage_im_out(102),
            data_im_out(4) => first_stage_im_out(134),
            data_im_out(5) => first_stage_im_out(166),
            data_im_out(6) => first_stage_im_out(198),
            data_im_out(7) => first_stage_im_out(230),
            data_im_out(8) => first_stage_im_out(262),
            data_im_out(9) => first_stage_im_out(294),
            data_im_out(10) => first_stage_im_out(326),
            data_im_out(11) => first_stage_im_out(358),
            data_im_out(12) => first_stage_im_out(390),
            data_im_out(13) => first_stage_im_out(422),
            data_im_out(14) => first_stage_im_out(454),
            data_im_out(15) => first_stage_im_out(486)
        );

    ULFFT_PT16_7 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(7),
            data_re_in(1) => data_re_in(39),
            data_re_in(2) => data_re_in(71),
            data_re_in(3) => data_re_in(103),
            data_re_in(4) => data_re_in(135),
            data_re_in(5) => data_re_in(167),
            data_re_in(6) => data_re_in(199),
            data_re_in(7) => data_re_in(231),
            data_re_in(8) => data_re_in(263),
            data_re_in(9) => data_re_in(295),
            data_re_in(10) => data_re_in(327),
            data_re_in(11) => data_re_in(359),
            data_re_in(12) => data_re_in(391),
            data_re_in(13) => data_re_in(423),
            data_re_in(14) => data_re_in(455),
            data_re_in(15) => data_re_in(487),
            data_im_in(0) => data_im_in(7),
            data_im_in(1) => data_im_in(39),
            data_im_in(2) => data_im_in(71),
            data_im_in(3) => data_im_in(103),
            data_im_in(4) => data_im_in(135),
            data_im_in(5) => data_im_in(167),
            data_im_in(6) => data_im_in(199),
            data_im_in(7) => data_im_in(231),
            data_im_in(8) => data_im_in(263),
            data_im_in(9) => data_im_in(295),
            data_im_in(10) => data_im_in(327),
            data_im_in(11) => data_im_in(359),
            data_im_in(12) => data_im_in(391),
            data_im_in(13) => data_im_in(423),
            data_im_in(14) => data_im_in(455),
            data_im_in(15) => data_im_in(487),
            data_re_out(0) => first_stage_re_out(7),
            data_re_out(1) => first_stage_re_out(39),
            data_re_out(2) => first_stage_re_out(71),
            data_re_out(3) => first_stage_re_out(103),
            data_re_out(4) => first_stage_re_out(135),
            data_re_out(5) => first_stage_re_out(167),
            data_re_out(6) => first_stage_re_out(199),
            data_re_out(7) => first_stage_re_out(231),
            data_re_out(8) => first_stage_re_out(263),
            data_re_out(9) => first_stage_re_out(295),
            data_re_out(10) => first_stage_re_out(327),
            data_re_out(11) => first_stage_re_out(359),
            data_re_out(12) => first_stage_re_out(391),
            data_re_out(13) => first_stage_re_out(423),
            data_re_out(14) => first_stage_re_out(455),
            data_re_out(15) => first_stage_re_out(487),
            data_im_out(0) => first_stage_im_out(7),
            data_im_out(1) => first_stage_im_out(39),
            data_im_out(2) => first_stage_im_out(71),
            data_im_out(3) => first_stage_im_out(103),
            data_im_out(4) => first_stage_im_out(135),
            data_im_out(5) => first_stage_im_out(167),
            data_im_out(6) => first_stage_im_out(199),
            data_im_out(7) => first_stage_im_out(231),
            data_im_out(8) => first_stage_im_out(263),
            data_im_out(9) => first_stage_im_out(295),
            data_im_out(10) => first_stage_im_out(327),
            data_im_out(11) => first_stage_im_out(359),
            data_im_out(12) => first_stage_im_out(391),
            data_im_out(13) => first_stage_im_out(423),
            data_im_out(14) => first_stage_im_out(455),
            data_im_out(15) => first_stage_im_out(487)
        );

    ULFFT_PT16_8 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(8),
            data_re_in(1) => data_re_in(40),
            data_re_in(2) => data_re_in(72),
            data_re_in(3) => data_re_in(104),
            data_re_in(4) => data_re_in(136),
            data_re_in(5) => data_re_in(168),
            data_re_in(6) => data_re_in(200),
            data_re_in(7) => data_re_in(232),
            data_re_in(8) => data_re_in(264),
            data_re_in(9) => data_re_in(296),
            data_re_in(10) => data_re_in(328),
            data_re_in(11) => data_re_in(360),
            data_re_in(12) => data_re_in(392),
            data_re_in(13) => data_re_in(424),
            data_re_in(14) => data_re_in(456),
            data_re_in(15) => data_re_in(488),
            data_im_in(0) => data_im_in(8),
            data_im_in(1) => data_im_in(40),
            data_im_in(2) => data_im_in(72),
            data_im_in(3) => data_im_in(104),
            data_im_in(4) => data_im_in(136),
            data_im_in(5) => data_im_in(168),
            data_im_in(6) => data_im_in(200),
            data_im_in(7) => data_im_in(232),
            data_im_in(8) => data_im_in(264),
            data_im_in(9) => data_im_in(296),
            data_im_in(10) => data_im_in(328),
            data_im_in(11) => data_im_in(360),
            data_im_in(12) => data_im_in(392),
            data_im_in(13) => data_im_in(424),
            data_im_in(14) => data_im_in(456),
            data_im_in(15) => data_im_in(488),
            data_re_out(0) => first_stage_re_out(8),
            data_re_out(1) => first_stage_re_out(40),
            data_re_out(2) => first_stage_re_out(72),
            data_re_out(3) => first_stage_re_out(104),
            data_re_out(4) => first_stage_re_out(136),
            data_re_out(5) => first_stage_re_out(168),
            data_re_out(6) => first_stage_re_out(200),
            data_re_out(7) => first_stage_re_out(232),
            data_re_out(8) => first_stage_re_out(264),
            data_re_out(9) => first_stage_re_out(296),
            data_re_out(10) => first_stage_re_out(328),
            data_re_out(11) => first_stage_re_out(360),
            data_re_out(12) => first_stage_re_out(392),
            data_re_out(13) => first_stage_re_out(424),
            data_re_out(14) => first_stage_re_out(456),
            data_re_out(15) => first_stage_re_out(488),
            data_im_out(0) => first_stage_im_out(8),
            data_im_out(1) => first_stage_im_out(40),
            data_im_out(2) => first_stage_im_out(72),
            data_im_out(3) => first_stage_im_out(104),
            data_im_out(4) => first_stage_im_out(136),
            data_im_out(5) => first_stage_im_out(168),
            data_im_out(6) => first_stage_im_out(200),
            data_im_out(7) => first_stage_im_out(232),
            data_im_out(8) => first_stage_im_out(264),
            data_im_out(9) => first_stage_im_out(296),
            data_im_out(10) => first_stage_im_out(328),
            data_im_out(11) => first_stage_im_out(360),
            data_im_out(12) => first_stage_im_out(392),
            data_im_out(13) => first_stage_im_out(424),
            data_im_out(14) => first_stage_im_out(456),
            data_im_out(15) => first_stage_im_out(488)
        );

    ULFFT_PT16_9 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(9),
            data_re_in(1) => data_re_in(41),
            data_re_in(2) => data_re_in(73),
            data_re_in(3) => data_re_in(105),
            data_re_in(4) => data_re_in(137),
            data_re_in(5) => data_re_in(169),
            data_re_in(6) => data_re_in(201),
            data_re_in(7) => data_re_in(233),
            data_re_in(8) => data_re_in(265),
            data_re_in(9) => data_re_in(297),
            data_re_in(10) => data_re_in(329),
            data_re_in(11) => data_re_in(361),
            data_re_in(12) => data_re_in(393),
            data_re_in(13) => data_re_in(425),
            data_re_in(14) => data_re_in(457),
            data_re_in(15) => data_re_in(489),
            data_im_in(0) => data_im_in(9),
            data_im_in(1) => data_im_in(41),
            data_im_in(2) => data_im_in(73),
            data_im_in(3) => data_im_in(105),
            data_im_in(4) => data_im_in(137),
            data_im_in(5) => data_im_in(169),
            data_im_in(6) => data_im_in(201),
            data_im_in(7) => data_im_in(233),
            data_im_in(8) => data_im_in(265),
            data_im_in(9) => data_im_in(297),
            data_im_in(10) => data_im_in(329),
            data_im_in(11) => data_im_in(361),
            data_im_in(12) => data_im_in(393),
            data_im_in(13) => data_im_in(425),
            data_im_in(14) => data_im_in(457),
            data_im_in(15) => data_im_in(489),
            data_re_out(0) => first_stage_re_out(9),
            data_re_out(1) => first_stage_re_out(41),
            data_re_out(2) => first_stage_re_out(73),
            data_re_out(3) => first_stage_re_out(105),
            data_re_out(4) => first_stage_re_out(137),
            data_re_out(5) => first_stage_re_out(169),
            data_re_out(6) => first_stage_re_out(201),
            data_re_out(7) => first_stage_re_out(233),
            data_re_out(8) => first_stage_re_out(265),
            data_re_out(9) => first_stage_re_out(297),
            data_re_out(10) => first_stage_re_out(329),
            data_re_out(11) => first_stage_re_out(361),
            data_re_out(12) => first_stage_re_out(393),
            data_re_out(13) => first_stage_re_out(425),
            data_re_out(14) => first_stage_re_out(457),
            data_re_out(15) => first_stage_re_out(489),
            data_im_out(0) => first_stage_im_out(9),
            data_im_out(1) => first_stage_im_out(41),
            data_im_out(2) => first_stage_im_out(73),
            data_im_out(3) => first_stage_im_out(105),
            data_im_out(4) => first_stage_im_out(137),
            data_im_out(5) => first_stage_im_out(169),
            data_im_out(6) => first_stage_im_out(201),
            data_im_out(7) => first_stage_im_out(233),
            data_im_out(8) => first_stage_im_out(265),
            data_im_out(9) => first_stage_im_out(297),
            data_im_out(10) => first_stage_im_out(329),
            data_im_out(11) => first_stage_im_out(361),
            data_im_out(12) => first_stage_im_out(393),
            data_im_out(13) => first_stage_im_out(425),
            data_im_out(14) => first_stage_im_out(457),
            data_im_out(15) => first_stage_im_out(489)
        );

    ULFFT_PT16_10 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(10),
            data_re_in(1) => data_re_in(42),
            data_re_in(2) => data_re_in(74),
            data_re_in(3) => data_re_in(106),
            data_re_in(4) => data_re_in(138),
            data_re_in(5) => data_re_in(170),
            data_re_in(6) => data_re_in(202),
            data_re_in(7) => data_re_in(234),
            data_re_in(8) => data_re_in(266),
            data_re_in(9) => data_re_in(298),
            data_re_in(10) => data_re_in(330),
            data_re_in(11) => data_re_in(362),
            data_re_in(12) => data_re_in(394),
            data_re_in(13) => data_re_in(426),
            data_re_in(14) => data_re_in(458),
            data_re_in(15) => data_re_in(490),
            data_im_in(0) => data_im_in(10),
            data_im_in(1) => data_im_in(42),
            data_im_in(2) => data_im_in(74),
            data_im_in(3) => data_im_in(106),
            data_im_in(4) => data_im_in(138),
            data_im_in(5) => data_im_in(170),
            data_im_in(6) => data_im_in(202),
            data_im_in(7) => data_im_in(234),
            data_im_in(8) => data_im_in(266),
            data_im_in(9) => data_im_in(298),
            data_im_in(10) => data_im_in(330),
            data_im_in(11) => data_im_in(362),
            data_im_in(12) => data_im_in(394),
            data_im_in(13) => data_im_in(426),
            data_im_in(14) => data_im_in(458),
            data_im_in(15) => data_im_in(490),
            data_re_out(0) => first_stage_re_out(10),
            data_re_out(1) => first_stage_re_out(42),
            data_re_out(2) => first_stage_re_out(74),
            data_re_out(3) => first_stage_re_out(106),
            data_re_out(4) => first_stage_re_out(138),
            data_re_out(5) => first_stage_re_out(170),
            data_re_out(6) => first_stage_re_out(202),
            data_re_out(7) => first_stage_re_out(234),
            data_re_out(8) => first_stage_re_out(266),
            data_re_out(9) => first_stage_re_out(298),
            data_re_out(10) => first_stage_re_out(330),
            data_re_out(11) => first_stage_re_out(362),
            data_re_out(12) => first_stage_re_out(394),
            data_re_out(13) => first_stage_re_out(426),
            data_re_out(14) => first_stage_re_out(458),
            data_re_out(15) => first_stage_re_out(490),
            data_im_out(0) => first_stage_im_out(10),
            data_im_out(1) => first_stage_im_out(42),
            data_im_out(2) => first_stage_im_out(74),
            data_im_out(3) => first_stage_im_out(106),
            data_im_out(4) => first_stage_im_out(138),
            data_im_out(5) => first_stage_im_out(170),
            data_im_out(6) => first_stage_im_out(202),
            data_im_out(7) => first_stage_im_out(234),
            data_im_out(8) => first_stage_im_out(266),
            data_im_out(9) => first_stage_im_out(298),
            data_im_out(10) => first_stage_im_out(330),
            data_im_out(11) => first_stage_im_out(362),
            data_im_out(12) => first_stage_im_out(394),
            data_im_out(13) => first_stage_im_out(426),
            data_im_out(14) => first_stage_im_out(458),
            data_im_out(15) => first_stage_im_out(490)
        );

    ULFFT_PT16_11 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(11),
            data_re_in(1) => data_re_in(43),
            data_re_in(2) => data_re_in(75),
            data_re_in(3) => data_re_in(107),
            data_re_in(4) => data_re_in(139),
            data_re_in(5) => data_re_in(171),
            data_re_in(6) => data_re_in(203),
            data_re_in(7) => data_re_in(235),
            data_re_in(8) => data_re_in(267),
            data_re_in(9) => data_re_in(299),
            data_re_in(10) => data_re_in(331),
            data_re_in(11) => data_re_in(363),
            data_re_in(12) => data_re_in(395),
            data_re_in(13) => data_re_in(427),
            data_re_in(14) => data_re_in(459),
            data_re_in(15) => data_re_in(491),
            data_im_in(0) => data_im_in(11),
            data_im_in(1) => data_im_in(43),
            data_im_in(2) => data_im_in(75),
            data_im_in(3) => data_im_in(107),
            data_im_in(4) => data_im_in(139),
            data_im_in(5) => data_im_in(171),
            data_im_in(6) => data_im_in(203),
            data_im_in(7) => data_im_in(235),
            data_im_in(8) => data_im_in(267),
            data_im_in(9) => data_im_in(299),
            data_im_in(10) => data_im_in(331),
            data_im_in(11) => data_im_in(363),
            data_im_in(12) => data_im_in(395),
            data_im_in(13) => data_im_in(427),
            data_im_in(14) => data_im_in(459),
            data_im_in(15) => data_im_in(491),
            data_re_out(0) => first_stage_re_out(11),
            data_re_out(1) => first_stage_re_out(43),
            data_re_out(2) => first_stage_re_out(75),
            data_re_out(3) => first_stage_re_out(107),
            data_re_out(4) => first_stage_re_out(139),
            data_re_out(5) => first_stage_re_out(171),
            data_re_out(6) => first_stage_re_out(203),
            data_re_out(7) => first_stage_re_out(235),
            data_re_out(8) => first_stage_re_out(267),
            data_re_out(9) => first_stage_re_out(299),
            data_re_out(10) => first_stage_re_out(331),
            data_re_out(11) => first_stage_re_out(363),
            data_re_out(12) => first_stage_re_out(395),
            data_re_out(13) => first_stage_re_out(427),
            data_re_out(14) => first_stage_re_out(459),
            data_re_out(15) => first_stage_re_out(491),
            data_im_out(0) => first_stage_im_out(11),
            data_im_out(1) => first_stage_im_out(43),
            data_im_out(2) => first_stage_im_out(75),
            data_im_out(3) => first_stage_im_out(107),
            data_im_out(4) => first_stage_im_out(139),
            data_im_out(5) => first_stage_im_out(171),
            data_im_out(6) => first_stage_im_out(203),
            data_im_out(7) => first_stage_im_out(235),
            data_im_out(8) => first_stage_im_out(267),
            data_im_out(9) => first_stage_im_out(299),
            data_im_out(10) => first_stage_im_out(331),
            data_im_out(11) => first_stage_im_out(363),
            data_im_out(12) => first_stage_im_out(395),
            data_im_out(13) => first_stage_im_out(427),
            data_im_out(14) => first_stage_im_out(459),
            data_im_out(15) => first_stage_im_out(491)
        );

    ULFFT_PT16_12 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(12),
            data_re_in(1) => data_re_in(44),
            data_re_in(2) => data_re_in(76),
            data_re_in(3) => data_re_in(108),
            data_re_in(4) => data_re_in(140),
            data_re_in(5) => data_re_in(172),
            data_re_in(6) => data_re_in(204),
            data_re_in(7) => data_re_in(236),
            data_re_in(8) => data_re_in(268),
            data_re_in(9) => data_re_in(300),
            data_re_in(10) => data_re_in(332),
            data_re_in(11) => data_re_in(364),
            data_re_in(12) => data_re_in(396),
            data_re_in(13) => data_re_in(428),
            data_re_in(14) => data_re_in(460),
            data_re_in(15) => data_re_in(492),
            data_im_in(0) => data_im_in(12),
            data_im_in(1) => data_im_in(44),
            data_im_in(2) => data_im_in(76),
            data_im_in(3) => data_im_in(108),
            data_im_in(4) => data_im_in(140),
            data_im_in(5) => data_im_in(172),
            data_im_in(6) => data_im_in(204),
            data_im_in(7) => data_im_in(236),
            data_im_in(8) => data_im_in(268),
            data_im_in(9) => data_im_in(300),
            data_im_in(10) => data_im_in(332),
            data_im_in(11) => data_im_in(364),
            data_im_in(12) => data_im_in(396),
            data_im_in(13) => data_im_in(428),
            data_im_in(14) => data_im_in(460),
            data_im_in(15) => data_im_in(492),
            data_re_out(0) => first_stage_re_out(12),
            data_re_out(1) => first_stage_re_out(44),
            data_re_out(2) => first_stage_re_out(76),
            data_re_out(3) => first_stage_re_out(108),
            data_re_out(4) => first_stage_re_out(140),
            data_re_out(5) => first_stage_re_out(172),
            data_re_out(6) => first_stage_re_out(204),
            data_re_out(7) => first_stage_re_out(236),
            data_re_out(8) => first_stage_re_out(268),
            data_re_out(9) => first_stage_re_out(300),
            data_re_out(10) => first_stage_re_out(332),
            data_re_out(11) => first_stage_re_out(364),
            data_re_out(12) => first_stage_re_out(396),
            data_re_out(13) => first_stage_re_out(428),
            data_re_out(14) => first_stage_re_out(460),
            data_re_out(15) => first_stage_re_out(492),
            data_im_out(0) => first_stage_im_out(12),
            data_im_out(1) => first_stage_im_out(44),
            data_im_out(2) => first_stage_im_out(76),
            data_im_out(3) => first_stage_im_out(108),
            data_im_out(4) => first_stage_im_out(140),
            data_im_out(5) => first_stage_im_out(172),
            data_im_out(6) => first_stage_im_out(204),
            data_im_out(7) => first_stage_im_out(236),
            data_im_out(8) => first_stage_im_out(268),
            data_im_out(9) => first_stage_im_out(300),
            data_im_out(10) => first_stage_im_out(332),
            data_im_out(11) => first_stage_im_out(364),
            data_im_out(12) => first_stage_im_out(396),
            data_im_out(13) => first_stage_im_out(428),
            data_im_out(14) => first_stage_im_out(460),
            data_im_out(15) => first_stage_im_out(492)
        );

    ULFFT_PT16_13 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(13),
            data_re_in(1) => data_re_in(45),
            data_re_in(2) => data_re_in(77),
            data_re_in(3) => data_re_in(109),
            data_re_in(4) => data_re_in(141),
            data_re_in(5) => data_re_in(173),
            data_re_in(6) => data_re_in(205),
            data_re_in(7) => data_re_in(237),
            data_re_in(8) => data_re_in(269),
            data_re_in(9) => data_re_in(301),
            data_re_in(10) => data_re_in(333),
            data_re_in(11) => data_re_in(365),
            data_re_in(12) => data_re_in(397),
            data_re_in(13) => data_re_in(429),
            data_re_in(14) => data_re_in(461),
            data_re_in(15) => data_re_in(493),
            data_im_in(0) => data_im_in(13),
            data_im_in(1) => data_im_in(45),
            data_im_in(2) => data_im_in(77),
            data_im_in(3) => data_im_in(109),
            data_im_in(4) => data_im_in(141),
            data_im_in(5) => data_im_in(173),
            data_im_in(6) => data_im_in(205),
            data_im_in(7) => data_im_in(237),
            data_im_in(8) => data_im_in(269),
            data_im_in(9) => data_im_in(301),
            data_im_in(10) => data_im_in(333),
            data_im_in(11) => data_im_in(365),
            data_im_in(12) => data_im_in(397),
            data_im_in(13) => data_im_in(429),
            data_im_in(14) => data_im_in(461),
            data_im_in(15) => data_im_in(493),
            data_re_out(0) => first_stage_re_out(13),
            data_re_out(1) => first_stage_re_out(45),
            data_re_out(2) => first_stage_re_out(77),
            data_re_out(3) => first_stage_re_out(109),
            data_re_out(4) => first_stage_re_out(141),
            data_re_out(5) => first_stage_re_out(173),
            data_re_out(6) => first_stage_re_out(205),
            data_re_out(7) => first_stage_re_out(237),
            data_re_out(8) => first_stage_re_out(269),
            data_re_out(9) => first_stage_re_out(301),
            data_re_out(10) => first_stage_re_out(333),
            data_re_out(11) => first_stage_re_out(365),
            data_re_out(12) => first_stage_re_out(397),
            data_re_out(13) => first_stage_re_out(429),
            data_re_out(14) => first_stage_re_out(461),
            data_re_out(15) => first_stage_re_out(493),
            data_im_out(0) => first_stage_im_out(13),
            data_im_out(1) => first_stage_im_out(45),
            data_im_out(2) => first_stage_im_out(77),
            data_im_out(3) => first_stage_im_out(109),
            data_im_out(4) => first_stage_im_out(141),
            data_im_out(5) => first_stage_im_out(173),
            data_im_out(6) => first_stage_im_out(205),
            data_im_out(7) => first_stage_im_out(237),
            data_im_out(8) => first_stage_im_out(269),
            data_im_out(9) => first_stage_im_out(301),
            data_im_out(10) => first_stage_im_out(333),
            data_im_out(11) => first_stage_im_out(365),
            data_im_out(12) => first_stage_im_out(397),
            data_im_out(13) => first_stage_im_out(429),
            data_im_out(14) => first_stage_im_out(461),
            data_im_out(15) => first_stage_im_out(493)
        );

    ULFFT_PT16_14 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(14),
            data_re_in(1) => data_re_in(46),
            data_re_in(2) => data_re_in(78),
            data_re_in(3) => data_re_in(110),
            data_re_in(4) => data_re_in(142),
            data_re_in(5) => data_re_in(174),
            data_re_in(6) => data_re_in(206),
            data_re_in(7) => data_re_in(238),
            data_re_in(8) => data_re_in(270),
            data_re_in(9) => data_re_in(302),
            data_re_in(10) => data_re_in(334),
            data_re_in(11) => data_re_in(366),
            data_re_in(12) => data_re_in(398),
            data_re_in(13) => data_re_in(430),
            data_re_in(14) => data_re_in(462),
            data_re_in(15) => data_re_in(494),
            data_im_in(0) => data_im_in(14),
            data_im_in(1) => data_im_in(46),
            data_im_in(2) => data_im_in(78),
            data_im_in(3) => data_im_in(110),
            data_im_in(4) => data_im_in(142),
            data_im_in(5) => data_im_in(174),
            data_im_in(6) => data_im_in(206),
            data_im_in(7) => data_im_in(238),
            data_im_in(8) => data_im_in(270),
            data_im_in(9) => data_im_in(302),
            data_im_in(10) => data_im_in(334),
            data_im_in(11) => data_im_in(366),
            data_im_in(12) => data_im_in(398),
            data_im_in(13) => data_im_in(430),
            data_im_in(14) => data_im_in(462),
            data_im_in(15) => data_im_in(494),
            data_re_out(0) => first_stage_re_out(14),
            data_re_out(1) => first_stage_re_out(46),
            data_re_out(2) => first_stage_re_out(78),
            data_re_out(3) => first_stage_re_out(110),
            data_re_out(4) => first_stage_re_out(142),
            data_re_out(5) => first_stage_re_out(174),
            data_re_out(6) => first_stage_re_out(206),
            data_re_out(7) => first_stage_re_out(238),
            data_re_out(8) => first_stage_re_out(270),
            data_re_out(9) => first_stage_re_out(302),
            data_re_out(10) => first_stage_re_out(334),
            data_re_out(11) => first_stage_re_out(366),
            data_re_out(12) => first_stage_re_out(398),
            data_re_out(13) => first_stage_re_out(430),
            data_re_out(14) => first_stage_re_out(462),
            data_re_out(15) => first_stage_re_out(494),
            data_im_out(0) => first_stage_im_out(14),
            data_im_out(1) => first_stage_im_out(46),
            data_im_out(2) => first_stage_im_out(78),
            data_im_out(3) => first_stage_im_out(110),
            data_im_out(4) => first_stage_im_out(142),
            data_im_out(5) => first_stage_im_out(174),
            data_im_out(6) => first_stage_im_out(206),
            data_im_out(7) => first_stage_im_out(238),
            data_im_out(8) => first_stage_im_out(270),
            data_im_out(9) => first_stage_im_out(302),
            data_im_out(10) => first_stage_im_out(334),
            data_im_out(11) => first_stage_im_out(366),
            data_im_out(12) => first_stage_im_out(398),
            data_im_out(13) => first_stage_im_out(430),
            data_im_out(14) => first_stage_im_out(462),
            data_im_out(15) => first_stage_im_out(494)
        );

    ULFFT_PT16_15 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(15),
            data_re_in(1) => data_re_in(47),
            data_re_in(2) => data_re_in(79),
            data_re_in(3) => data_re_in(111),
            data_re_in(4) => data_re_in(143),
            data_re_in(5) => data_re_in(175),
            data_re_in(6) => data_re_in(207),
            data_re_in(7) => data_re_in(239),
            data_re_in(8) => data_re_in(271),
            data_re_in(9) => data_re_in(303),
            data_re_in(10) => data_re_in(335),
            data_re_in(11) => data_re_in(367),
            data_re_in(12) => data_re_in(399),
            data_re_in(13) => data_re_in(431),
            data_re_in(14) => data_re_in(463),
            data_re_in(15) => data_re_in(495),
            data_im_in(0) => data_im_in(15),
            data_im_in(1) => data_im_in(47),
            data_im_in(2) => data_im_in(79),
            data_im_in(3) => data_im_in(111),
            data_im_in(4) => data_im_in(143),
            data_im_in(5) => data_im_in(175),
            data_im_in(6) => data_im_in(207),
            data_im_in(7) => data_im_in(239),
            data_im_in(8) => data_im_in(271),
            data_im_in(9) => data_im_in(303),
            data_im_in(10) => data_im_in(335),
            data_im_in(11) => data_im_in(367),
            data_im_in(12) => data_im_in(399),
            data_im_in(13) => data_im_in(431),
            data_im_in(14) => data_im_in(463),
            data_im_in(15) => data_im_in(495),
            data_re_out(0) => first_stage_re_out(15),
            data_re_out(1) => first_stage_re_out(47),
            data_re_out(2) => first_stage_re_out(79),
            data_re_out(3) => first_stage_re_out(111),
            data_re_out(4) => first_stage_re_out(143),
            data_re_out(5) => first_stage_re_out(175),
            data_re_out(6) => first_stage_re_out(207),
            data_re_out(7) => first_stage_re_out(239),
            data_re_out(8) => first_stage_re_out(271),
            data_re_out(9) => first_stage_re_out(303),
            data_re_out(10) => first_stage_re_out(335),
            data_re_out(11) => first_stage_re_out(367),
            data_re_out(12) => first_stage_re_out(399),
            data_re_out(13) => first_stage_re_out(431),
            data_re_out(14) => first_stage_re_out(463),
            data_re_out(15) => first_stage_re_out(495),
            data_im_out(0) => first_stage_im_out(15),
            data_im_out(1) => first_stage_im_out(47),
            data_im_out(2) => first_stage_im_out(79),
            data_im_out(3) => first_stage_im_out(111),
            data_im_out(4) => first_stage_im_out(143),
            data_im_out(5) => first_stage_im_out(175),
            data_im_out(6) => first_stage_im_out(207),
            data_im_out(7) => first_stage_im_out(239),
            data_im_out(8) => first_stage_im_out(271),
            data_im_out(9) => first_stage_im_out(303),
            data_im_out(10) => first_stage_im_out(335),
            data_im_out(11) => first_stage_im_out(367),
            data_im_out(12) => first_stage_im_out(399),
            data_im_out(13) => first_stage_im_out(431),
            data_im_out(14) => first_stage_im_out(463),
            data_im_out(15) => first_stage_im_out(495)
        );

    ULFFT_PT16_16 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(16),
            data_re_in(1) => data_re_in(48),
            data_re_in(2) => data_re_in(80),
            data_re_in(3) => data_re_in(112),
            data_re_in(4) => data_re_in(144),
            data_re_in(5) => data_re_in(176),
            data_re_in(6) => data_re_in(208),
            data_re_in(7) => data_re_in(240),
            data_re_in(8) => data_re_in(272),
            data_re_in(9) => data_re_in(304),
            data_re_in(10) => data_re_in(336),
            data_re_in(11) => data_re_in(368),
            data_re_in(12) => data_re_in(400),
            data_re_in(13) => data_re_in(432),
            data_re_in(14) => data_re_in(464),
            data_re_in(15) => data_re_in(496),
            data_im_in(0) => data_im_in(16),
            data_im_in(1) => data_im_in(48),
            data_im_in(2) => data_im_in(80),
            data_im_in(3) => data_im_in(112),
            data_im_in(4) => data_im_in(144),
            data_im_in(5) => data_im_in(176),
            data_im_in(6) => data_im_in(208),
            data_im_in(7) => data_im_in(240),
            data_im_in(8) => data_im_in(272),
            data_im_in(9) => data_im_in(304),
            data_im_in(10) => data_im_in(336),
            data_im_in(11) => data_im_in(368),
            data_im_in(12) => data_im_in(400),
            data_im_in(13) => data_im_in(432),
            data_im_in(14) => data_im_in(464),
            data_im_in(15) => data_im_in(496),
            data_re_out(0) => first_stage_re_out(16),
            data_re_out(1) => first_stage_re_out(48),
            data_re_out(2) => first_stage_re_out(80),
            data_re_out(3) => first_stage_re_out(112),
            data_re_out(4) => first_stage_re_out(144),
            data_re_out(5) => first_stage_re_out(176),
            data_re_out(6) => first_stage_re_out(208),
            data_re_out(7) => first_stage_re_out(240),
            data_re_out(8) => first_stage_re_out(272),
            data_re_out(9) => first_stage_re_out(304),
            data_re_out(10) => first_stage_re_out(336),
            data_re_out(11) => first_stage_re_out(368),
            data_re_out(12) => first_stage_re_out(400),
            data_re_out(13) => first_stage_re_out(432),
            data_re_out(14) => first_stage_re_out(464),
            data_re_out(15) => first_stage_re_out(496),
            data_im_out(0) => first_stage_im_out(16),
            data_im_out(1) => first_stage_im_out(48),
            data_im_out(2) => first_stage_im_out(80),
            data_im_out(3) => first_stage_im_out(112),
            data_im_out(4) => first_stage_im_out(144),
            data_im_out(5) => first_stage_im_out(176),
            data_im_out(6) => first_stage_im_out(208),
            data_im_out(7) => first_stage_im_out(240),
            data_im_out(8) => first_stage_im_out(272),
            data_im_out(9) => first_stage_im_out(304),
            data_im_out(10) => first_stage_im_out(336),
            data_im_out(11) => first_stage_im_out(368),
            data_im_out(12) => first_stage_im_out(400),
            data_im_out(13) => first_stage_im_out(432),
            data_im_out(14) => first_stage_im_out(464),
            data_im_out(15) => first_stage_im_out(496)
        );

    ULFFT_PT16_17 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(17),
            data_re_in(1) => data_re_in(49),
            data_re_in(2) => data_re_in(81),
            data_re_in(3) => data_re_in(113),
            data_re_in(4) => data_re_in(145),
            data_re_in(5) => data_re_in(177),
            data_re_in(6) => data_re_in(209),
            data_re_in(7) => data_re_in(241),
            data_re_in(8) => data_re_in(273),
            data_re_in(9) => data_re_in(305),
            data_re_in(10) => data_re_in(337),
            data_re_in(11) => data_re_in(369),
            data_re_in(12) => data_re_in(401),
            data_re_in(13) => data_re_in(433),
            data_re_in(14) => data_re_in(465),
            data_re_in(15) => data_re_in(497),
            data_im_in(0) => data_im_in(17),
            data_im_in(1) => data_im_in(49),
            data_im_in(2) => data_im_in(81),
            data_im_in(3) => data_im_in(113),
            data_im_in(4) => data_im_in(145),
            data_im_in(5) => data_im_in(177),
            data_im_in(6) => data_im_in(209),
            data_im_in(7) => data_im_in(241),
            data_im_in(8) => data_im_in(273),
            data_im_in(9) => data_im_in(305),
            data_im_in(10) => data_im_in(337),
            data_im_in(11) => data_im_in(369),
            data_im_in(12) => data_im_in(401),
            data_im_in(13) => data_im_in(433),
            data_im_in(14) => data_im_in(465),
            data_im_in(15) => data_im_in(497),
            data_re_out(0) => first_stage_re_out(17),
            data_re_out(1) => first_stage_re_out(49),
            data_re_out(2) => first_stage_re_out(81),
            data_re_out(3) => first_stage_re_out(113),
            data_re_out(4) => first_stage_re_out(145),
            data_re_out(5) => first_stage_re_out(177),
            data_re_out(6) => first_stage_re_out(209),
            data_re_out(7) => first_stage_re_out(241),
            data_re_out(8) => first_stage_re_out(273),
            data_re_out(9) => first_stage_re_out(305),
            data_re_out(10) => first_stage_re_out(337),
            data_re_out(11) => first_stage_re_out(369),
            data_re_out(12) => first_stage_re_out(401),
            data_re_out(13) => first_stage_re_out(433),
            data_re_out(14) => first_stage_re_out(465),
            data_re_out(15) => first_stage_re_out(497),
            data_im_out(0) => first_stage_im_out(17),
            data_im_out(1) => first_stage_im_out(49),
            data_im_out(2) => first_stage_im_out(81),
            data_im_out(3) => first_stage_im_out(113),
            data_im_out(4) => first_stage_im_out(145),
            data_im_out(5) => first_stage_im_out(177),
            data_im_out(6) => first_stage_im_out(209),
            data_im_out(7) => first_stage_im_out(241),
            data_im_out(8) => first_stage_im_out(273),
            data_im_out(9) => first_stage_im_out(305),
            data_im_out(10) => first_stage_im_out(337),
            data_im_out(11) => first_stage_im_out(369),
            data_im_out(12) => first_stage_im_out(401),
            data_im_out(13) => first_stage_im_out(433),
            data_im_out(14) => first_stage_im_out(465),
            data_im_out(15) => first_stage_im_out(497)
        );

    ULFFT_PT16_18 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(18),
            data_re_in(1) => data_re_in(50),
            data_re_in(2) => data_re_in(82),
            data_re_in(3) => data_re_in(114),
            data_re_in(4) => data_re_in(146),
            data_re_in(5) => data_re_in(178),
            data_re_in(6) => data_re_in(210),
            data_re_in(7) => data_re_in(242),
            data_re_in(8) => data_re_in(274),
            data_re_in(9) => data_re_in(306),
            data_re_in(10) => data_re_in(338),
            data_re_in(11) => data_re_in(370),
            data_re_in(12) => data_re_in(402),
            data_re_in(13) => data_re_in(434),
            data_re_in(14) => data_re_in(466),
            data_re_in(15) => data_re_in(498),
            data_im_in(0) => data_im_in(18),
            data_im_in(1) => data_im_in(50),
            data_im_in(2) => data_im_in(82),
            data_im_in(3) => data_im_in(114),
            data_im_in(4) => data_im_in(146),
            data_im_in(5) => data_im_in(178),
            data_im_in(6) => data_im_in(210),
            data_im_in(7) => data_im_in(242),
            data_im_in(8) => data_im_in(274),
            data_im_in(9) => data_im_in(306),
            data_im_in(10) => data_im_in(338),
            data_im_in(11) => data_im_in(370),
            data_im_in(12) => data_im_in(402),
            data_im_in(13) => data_im_in(434),
            data_im_in(14) => data_im_in(466),
            data_im_in(15) => data_im_in(498),
            data_re_out(0) => first_stage_re_out(18),
            data_re_out(1) => first_stage_re_out(50),
            data_re_out(2) => first_stage_re_out(82),
            data_re_out(3) => first_stage_re_out(114),
            data_re_out(4) => first_stage_re_out(146),
            data_re_out(5) => first_stage_re_out(178),
            data_re_out(6) => first_stage_re_out(210),
            data_re_out(7) => first_stage_re_out(242),
            data_re_out(8) => first_stage_re_out(274),
            data_re_out(9) => first_stage_re_out(306),
            data_re_out(10) => first_stage_re_out(338),
            data_re_out(11) => first_stage_re_out(370),
            data_re_out(12) => first_stage_re_out(402),
            data_re_out(13) => first_stage_re_out(434),
            data_re_out(14) => first_stage_re_out(466),
            data_re_out(15) => first_stage_re_out(498),
            data_im_out(0) => first_stage_im_out(18),
            data_im_out(1) => first_stage_im_out(50),
            data_im_out(2) => first_stage_im_out(82),
            data_im_out(3) => first_stage_im_out(114),
            data_im_out(4) => first_stage_im_out(146),
            data_im_out(5) => first_stage_im_out(178),
            data_im_out(6) => first_stage_im_out(210),
            data_im_out(7) => first_stage_im_out(242),
            data_im_out(8) => first_stage_im_out(274),
            data_im_out(9) => first_stage_im_out(306),
            data_im_out(10) => first_stage_im_out(338),
            data_im_out(11) => first_stage_im_out(370),
            data_im_out(12) => first_stage_im_out(402),
            data_im_out(13) => first_stage_im_out(434),
            data_im_out(14) => first_stage_im_out(466),
            data_im_out(15) => first_stage_im_out(498)
        );

    ULFFT_PT16_19 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(19),
            data_re_in(1) => data_re_in(51),
            data_re_in(2) => data_re_in(83),
            data_re_in(3) => data_re_in(115),
            data_re_in(4) => data_re_in(147),
            data_re_in(5) => data_re_in(179),
            data_re_in(6) => data_re_in(211),
            data_re_in(7) => data_re_in(243),
            data_re_in(8) => data_re_in(275),
            data_re_in(9) => data_re_in(307),
            data_re_in(10) => data_re_in(339),
            data_re_in(11) => data_re_in(371),
            data_re_in(12) => data_re_in(403),
            data_re_in(13) => data_re_in(435),
            data_re_in(14) => data_re_in(467),
            data_re_in(15) => data_re_in(499),
            data_im_in(0) => data_im_in(19),
            data_im_in(1) => data_im_in(51),
            data_im_in(2) => data_im_in(83),
            data_im_in(3) => data_im_in(115),
            data_im_in(4) => data_im_in(147),
            data_im_in(5) => data_im_in(179),
            data_im_in(6) => data_im_in(211),
            data_im_in(7) => data_im_in(243),
            data_im_in(8) => data_im_in(275),
            data_im_in(9) => data_im_in(307),
            data_im_in(10) => data_im_in(339),
            data_im_in(11) => data_im_in(371),
            data_im_in(12) => data_im_in(403),
            data_im_in(13) => data_im_in(435),
            data_im_in(14) => data_im_in(467),
            data_im_in(15) => data_im_in(499),
            data_re_out(0) => first_stage_re_out(19),
            data_re_out(1) => first_stage_re_out(51),
            data_re_out(2) => first_stage_re_out(83),
            data_re_out(3) => first_stage_re_out(115),
            data_re_out(4) => first_stage_re_out(147),
            data_re_out(5) => first_stage_re_out(179),
            data_re_out(6) => first_stage_re_out(211),
            data_re_out(7) => first_stage_re_out(243),
            data_re_out(8) => first_stage_re_out(275),
            data_re_out(9) => first_stage_re_out(307),
            data_re_out(10) => first_stage_re_out(339),
            data_re_out(11) => first_stage_re_out(371),
            data_re_out(12) => first_stage_re_out(403),
            data_re_out(13) => first_stage_re_out(435),
            data_re_out(14) => first_stage_re_out(467),
            data_re_out(15) => first_stage_re_out(499),
            data_im_out(0) => first_stage_im_out(19),
            data_im_out(1) => first_stage_im_out(51),
            data_im_out(2) => first_stage_im_out(83),
            data_im_out(3) => first_stage_im_out(115),
            data_im_out(4) => first_stage_im_out(147),
            data_im_out(5) => first_stage_im_out(179),
            data_im_out(6) => first_stage_im_out(211),
            data_im_out(7) => first_stage_im_out(243),
            data_im_out(8) => first_stage_im_out(275),
            data_im_out(9) => first_stage_im_out(307),
            data_im_out(10) => first_stage_im_out(339),
            data_im_out(11) => first_stage_im_out(371),
            data_im_out(12) => first_stage_im_out(403),
            data_im_out(13) => first_stage_im_out(435),
            data_im_out(14) => first_stage_im_out(467),
            data_im_out(15) => first_stage_im_out(499)
        );

    ULFFT_PT16_20 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(20),
            data_re_in(1) => data_re_in(52),
            data_re_in(2) => data_re_in(84),
            data_re_in(3) => data_re_in(116),
            data_re_in(4) => data_re_in(148),
            data_re_in(5) => data_re_in(180),
            data_re_in(6) => data_re_in(212),
            data_re_in(7) => data_re_in(244),
            data_re_in(8) => data_re_in(276),
            data_re_in(9) => data_re_in(308),
            data_re_in(10) => data_re_in(340),
            data_re_in(11) => data_re_in(372),
            data_re_in(12) => data_re_in(404),
            data_re_in(13) => data_re_in(436),
            data_re_in(14) => data_re_in(468),
            data_re_in(15) => data_re_in(500),
            data_im_in(0) => data_im_in(20),
            data_im_in(1) => data_im_in(52),
            data_im_in(2) => data_im_in(84),
            data_im_in(3) => data_im_in(116),
            data_im_in(4) => data_im_in(148),
            data_im_in(5) => data_im_in(180),
            data_im_in(6) => data_im_in(212),
            data_im_in(7) => data_im_in(244),
            data_im_in(8) => data_im_in(276),
            data_im_in(9) => data_im_in(308),
            data_im_in(10) => data_im_in(340),
            data_im_in(11) => data_im_in(372),
            data_im_in(12) => data_im_in(404),
            data_im_in(13) => data_im_in(436),
            data_im_in(14) => data_im_in(468),
            data_im_in(15) => data_im_in(500),
            data_re_out(0) => first_stage_re_out(20),
            data_re_out(1) => first_stage_re_out(52),
            data_re_out(2) => first_stage_re_out(84),
            data_re_out(3) => first_stage_re_out(116),
            data_re_out(4) => first_stage_re_out(148),
            data_re_out(5) => first_stage_re_out(180),
            data_re_out(6) => first_stage_re_out(212),
            data_re_out(7) => first_stage_re_out(244),
            data_re_out(8) => first_stage_re_out(276),
            data_re_out(9) => first_stage_re_out(308),
            data_re_out(10) => first_stage_re_out(340),
            data_re_out(11) => first_stage_re_out(372),
            data_re_out(12) => first_stage_re_out(404),
            data_re_out(13) => first_stage_re_out(436),
            data_re_out(14) => first_stage_re_out(468),
            data_re_out(15) => first_stage_re_out(500),
            data_im_out(0) => first_stage_im_out(20),
            data_im_out(1) => first_stage_im_out(52),
            data_im_out(2) => first_stage_im_out(84),
            data_im_out(3) => first_stage_im_out(116),
            data_im_out(4) => first_stage_im_out(148),
            data_im_out(5) => first_stage_im_out(180),
            data_im_out(6) => first_stage_im_out(212),
            data_im_out(7) => first_stage_im_out(244),
            data_im_out(8) => first_stage_im_out(276),
            data_im_out(9) => first_stage_im_out(308),
            data_im_out(10) => first_stage_im_out(340),
            data_im_out(11) => first_stage_im_out(372),
            data_im_out(12) => first_stage_im_out(404),
            data_im_out(13) => first_stage_im_out(436),
            data_im_out(14) => first_stage_im_out(468),
            data_im_out(15) => first_stage_im_out(500)
        );

    ULFFT_PT16_21 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(21),
            data_re_in(1) => data_re_in(53),
            data_re_in(2) => data_re_in(85),
            data_re_in(3) => data_re_in(117),
            data_re_in(4) => data_re_in(149),
            data_re_in(5) => data_re_in(181),
            data_re_in(6) => data_re_in(213),
            data_re_in(7) => data_re_in(245),
            data_re_in(8) => data_re_in(277),
            data_re_in(9) => data_re_in(309),
            data_re_in(10) => data_re_in(341),
            data_re_in(11) => data_re_in(373),
            data_re_in(12) => data_re_in(405),
            data_re_in(13) => data_re_in(437),
            data_re_in(14) => data_re_in(469),
            data_re_in(15) => data_re_in(501),
            data_im_in(0) => data_im_in(21),
            data_im_in(1) => data_im_in(53),
            data_im_in(2) => data_im_in(85),
            data_im_in(3) => data_im_in(117),
            data_im_in(4) => data_im_in(149),
            data_im_in(5) => data_im_in(181),
            data_im_in(6) => data_im_in(213),
            data_im_in(7) => data_im_in(245),
            data_im_in(8) => data_im_in(277),
            data_im_in(9) => data_im_in(309),
            data_im_in(10) => data_im_in(341),
            data_im_in(11) => data_im_in(373),
            data_im_in(12) => data_im_in(405),
            data_im_in(13) => data_im_in(437),
            data_im_in(14) => data_im_in(469),
            data_im_in(15) => data_im_in(501),
            data_re_out(0) => first_stage_re_out(21),
            data_re_out(1) => first_stage_re_out(53),
            data_re_out(2) => first_stage_re_out(85),
            data_re_out(3) => first_stage_re_out(117),
            data_re_out(4) => first_stage_re_out(149),
            data_re_out(5) => first_stage_re_out(181),
            data_re_out(6) => first_stage_re_out(213),
            data_re_out(7) => first_stage_re_out(245),
            data_re_out(8) => first_stage_re_out(277),
            data_re_out(9) => first_stage_re_out(309),
            data_re_out(10) => first_stage_re_out(341),
            data_re_out(11) => first_stage_re_out(373),
            data_re_out(12) => first_stage_re_out(405),
            data_re_out(13) => first_stage_re_out(437),
            data_re_out(14) => first_stage_re_out(469),
            data_re_out(15) => first_stage_re_out(501),
            data_im_out(0) => first_stage_im_out(21),
            data_im_out(1) => first_stage_im_out(53),
            data_im_out(2) => first_stage_im_out(85),
            data_im_out(3) => first_stage_im_out(117),
            data_im_out(4) => first_stage_im_out(149),
            data_im_out(5) => first_stage_im_out(181),
            data_im_out(6) => first_stage_im_out(213),
            data_im_out(7) => first_stage_im_out(245),
            data_im_out(8) => first_stage_im_out(277),
            data_im_out(9) => first_stage_im_out(309),
            data_im_out(10) => first_stage_im_out(341),
            data_im_out(11) => first_stage_im_out(373),
            data_im_out(12) => first_stage_im_out(405),
            data_im_out(13) => first_stage_im_out(437),
            data_im_out(14) => first_stage_im_out(469),
            data_im_out(15) => first_stage_im_out(501)
        );

    ULFFT_PT16_22 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(22),
            data_re_in(1) => data_re_in(54),
            data_re_in(2) => data_re_in(86),
            data_re_in(3) => data_re_in(118),
            data_re_in(4) => data_re_in(150),
            data_re_in(5) => data_re_in(182),
            data_re_in(6) => data_re_in(214),
            data_re_in(7) => data_re_in(246),
            data_re_in(8) => data_re_in(278),
            data_re_in(9) => data_re_in(310),
            data_re_in(10) => data_re_in(342),
            data_re_in(11) => data_re_in(374),
            data_re_in(12) => data_re_in(406),
            data_re_in(13) => data_re_in(438),
            data_re_in(14) => data_re_in(470),
            data_re_in(15) => data_re_in(502),
            data_im_in(0) => data_im_in(22),
            data_im_in(1) => data_im_in(54),
            data_im_in(2) => data_im_in(86),
            data_im_in(3) => data_im_in(118),
            data_im_in(4) => data_im_in(150),
            data_im_in(5) => data_im_in(182),
            data_im_in(6) => data_im_in(214),
            data_im_in(7) => data_im_in(246),
            data_im_in(8) => data_im_in(278),
            data_im_in(9) => data_im_in(310),
            data_im_in(10) => data_im_in(342),
            data_im_in(11) => data_im_in(374),
            data_im_in(12) => data_im_in(406),
            data_im_in(13) => data_im_in(438),
            data_im_in(14) => data_im_in(470),
            data_im_in(15) => data_im_in(502),
            data_re_out(0) => first_stage_re_out(22),
            data_re_out(1) => first_stage_re_out(54),
            data_re_out(2) => first_stage_re_out(86),
            data_re_out(3) => first_stage_re_out(118),
            data_re_out(4) => first_stage_re_out(150),
            data_re_out(5) => first_stage_re_out(182),
            data_re_out(6) => first_stage_re_out(214),
            data_re_out(7) => first_stage_re_out(246),
            data_re_out(8) => first_stage_re_out(278),
            data_re_out(9) => first_stage_re_out(310),
            data_re_out(10) => first_stage_re_out(342),
            data_re_out(11) => first_stage_re_out(374),
            data_re_out(12) => first_stage_re_out(406),
            data_re_out(13) => first_stage_re_out(438),
            data_re_out(14) => first_stage_re_out(470),
            data_re_out(15) => first_stage_re_out(502),
            data_im_out(0) => first_stage_im_out(22),
            data_im_out(1) => first_stage_im_out(54),
            data_im_out(2) => first_stage_im_out(86),
            data_im_out(3) => first_stage_im_out(118),
            data_im_out(4) => first_stage_im_out(150),
            data_im_out(5) => first_stage_im_out(182),
            data_im_out(6) => first_stage_im_out(214),
            data_im_out(7) => first_stage_im_out(246),
            data_im_out(8) => first_stage_im_out(278),
            data_im_out(9) => first_stage_im_out(310),
            data_im_out(10) => first_stage_im_out(342),
            data_im_out(11) => first_stage_im_out(374),
            data_im_out(12) => first_stage_im_out(406),
            data_im_out(13) => first_stage_im_out(438),
            data_im_out(14) => first_stage_im_out(470),
            data_im_out(15) => first_stage_im_out(502)
        );

    ULFFT_PT16_23 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(23),
            data_re_in(1) => data_re_in(55),
            data_re_in(2) => data_re_in(87),
            data_re_in(3) => data_re_in(119),
            data_re_in(4) => data_re_in(151),
            data_re_in(5) => data_re_in(183),
            data_re_in(6) => data_re_in(215),
            data_re_in(7) => data_re_in(247),
            data_re_in(8) => data_re_in(279),
            data_re_in(9) => data_re_in(311),
            data_re_in(10) => data_re_in(343),
            data_re_in(11) => data_re_in(375),
            data_re_in(12) => data_re_in(407),
            data_re_in(13) => data_re_in(439),
            data_re_in(14) => data_re_in(471),
            data_re_in(15) => data_re_in(503),
            data_im_in(0) => data_im_in(23),
            data_im_in(1) => data_im_in(55),
            data_im_in(2) => data_im_in(87),
            data_im_in(3) => data_im_in(119),
            data_im_in(4) => data_im_in(151),
            data_im_in(5) => data_im_in(183),
            data_im_in(6) => data_im_in(215),
            data_im_in(7) => data_im_in(247),
            data_im_in(8) => data_im_in(279),
            data_im_in(9) => data_im_in(311),
            data_im_in(10) => data_im_in(343),
            data_im_in(11) => data_im_in(375),
            data_im_in(12) => data_im_in(407),
            data_im_in(13) => data_im_in(439),
            data_im_in(14) => data_im_in(471),
            data_im_in(15) => data_im_in(503),
            data_re_out(0) => first_stage_re_out(23),
            data_re_out(1) => first_stage_re_out(55),
            data_re_out(2) => first_stage_re_out(87),
            data_re_out(3) => first_stage_re_out(119),
            data_re_out(4) => first_stage_re_out(151),
            data_re_out(5) => first_stage_re_out(183),
            data_re_out(6) => first_stage_re_out(215),
            data_re_out(7) => first_stage_re_out(247),
            data_re_out(8) => first_stage_re_out(279),
            data_re_out(9) => first_stage_re_out(311),
            data_re_out(10) => first_stage_re_out(343),
            data_re_out(11) => first_stage_re_out(375),
            data_re_out(12) => first_stage_re_out(407),
            data_re_out(13) => first_stage_re_out(439),
            data_re_out(14) => first_stage_re_out(471),
            data_re_out(15) => first_stage_re_out(503),
            data_im_out(0) => first_stage_im_out(23),
            data_im_out(1) => first_stage_im_out(55),
            data_im_out(2) => first_stage_im_out(87),
            data_im_out(3) => first_stage_im_out(119),
            data_im_out(4) => first_stage_im_out(151),
            data_im_out(5) => first_stage_im_out(183),
            data_im_out(6) => first_stage_im_out(215),
            data_im_out(7) => first_stage_im_out(247),
            data_im_out(8) => first_stage_im_out(279),
            data_im_out(9) => first_stage_im_out(311),
            data_im_out(10) => first_stage_im_out(343),
            data_im_out(11) => first_stage_im_out(375),
            data_im_out(12) => first_stage_im_out(407),
            data_im_out(13) => first_stage_im_out(439),
            data_im_out(14) => first_stage_im_out(471),
            data_im_out(15) => first_stage_im_out(503)
        );

    ULFFT_PT16_24 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(24),
            data_re_in(1) => data_re_in(56),
            data_re_in(2) => data_re_in(88),
            data_re_in(3) => data_re_in(120),
            data_re_in(4) => data_re_in(152),
            data_re_in(5) => data_re_in(184),
            data_re_in(6) => data_re_in(216),
            data_re_in(7) => data_re_in(248),
            data_re_in(8) => data_re_in(280),
            data_re_in(9) => data_re_in(312),
            data_re_in(10) => data_re_in(344),
            data_re_in(11) => data_re_in(376),
            data_re_in(12) => data_re_in(408),
            data_re_in(13) => data_re_in(440),
            data_re_in(14) => data_re_in(472),
            data_re_in(15) => data_re_in(504),
            data_im_in(0) => data_im_in(24),
            data_im_in(1) => data_im_in(56),
            data_im_in(2) => data_im_in(88),
            data_im_in(3) => data_im_in(120),
            data_im_in(4) => data_im_in(152),
            data_im_in(5) => data_im_in(184),
            data_im_in(6) => data_im_in(216),
            data_im_in(7) => data_im_in(248),
            data_im_in(8) => data_im_in(280),
            data_im_in(9) => data_im_in(312),
            data_im_in(10) => data_im_in(344),
            data_im_in(11) => data_im_in(376),
            data_im_in(12) => data_im_in(408),
            data_im_in(13) => data_im_in(440),
            data_im_in(14) => data_im_in(472),
            data_im_in(15) => data_im_in(504),
            data_re_out(0) => first_stage_re_out(24),
            data_re_out(1) => first_stage_re_out(56),
            data_re_out(2) => first_stage_re_out(88),
            data_re_out(3) => first_stage_re_out(120),
            data_re_out(4) => first_stage_re_out(152),
            data_re_out(5) => first_stage_re_out(184),
            data_re_out(6) => first_stage_re_out(216),
            data_re_out(7) => first_stage_re_out(248),
            data_re_out(8) => first_stage_re_out(280),
            data_re_out(9) => first_stage_re_out(312),
            data_re_out(10) => first_stage_re_out(344),
            data_re_out(11) => first_stage_re_out(376),
            data_re_out(12) => first_stage_re_out(408),
            data_re_out(13) => first_stage_re_out(440),
            data_re_out(14) => first_stage_re_out(472),
            data_re_out(15) => first_stage_re_out(504),
            data_im_out(0) => first_stage_im_out(24),
            data_im_out(1) => first_stage_im_out(56),
            data_im_out(2) => first_stage_im_out(88),
            data_im_out(3) => first_stage_im_out(120),
            data_im_out(4) => first_stage_im_out(152),
            data_im_out(5) => first_stage_im_out(184),
            data_im_out(6) => first_stage_im_out(216),
            data_im_out(7) => first_stage_im_out(248),
            data_im_out(8) => first_stage_im_out(280),
            data_im_out(9) => first_stage_im_out(312),
            data_im_out(10) => first_stage_im_out(344),
            data_im_out(11) => first_stage_im_out(376),
            data_im_out(12) => first_stage_im_out(408),
            data_im_out(13) => first_stage_im_out(440),
            data_im_out(14) => first_stage_im_out(472),
            data_im_out(15) => first_stage_im_out(504)
        );

    ULFFT_PT16_25 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(25),
            data_re_in(1) => data_re_in(57),
            data_re_in(2) => data_re_in(89),
            data_re_in(3) => data_re_in(121),
            data_re_in(4) => data_re_in(153),
            data_re_in(5) => data_re_in(185),
            data_re_in(6) => data_re_in(217),
            data_re_in(7) => data_re_in(249),
            data_re_in(8) => data_re_in(281),
            data_re_in(9) => data_re_in(313),
            data_re_in(10) => data_re_in(345),
            data_re_in(11) => data_re_in(377),
            data_re_in(12) => data_re_in(409),
            data_re_in(13) => data_re_in(441),
            data_re_in(14) => data_re_in(473),
            data_re_in(15) => data_re_in(505),
            data_im_in(0) => data_im_in(25),
            data_im_in(1) => data_im_in(57),
            data_im_in(2) => data_im_in(89),
            data_im_in(3) => data_im_in(121),
            data_im_in(4) => data_im_in(153),
            data_im_in(5) => data_im_in(185),
            data_im_in(6) => data_im_in(217),
            data_im_in(7) => data_im_in(249),
            data_im_in(8) => data_im_in(281),
            data_im_in(9) => data_im_in(313),
            data_im_in(10) => data_im_in(345),
            data_im_in(11) => data_im_in(377),
            data_im_in(12) => data_im_in(409),
            data_im_in(13) => data_im_in(441),
            data_im_in(14) => data_im_in(473),
            data_im_in(15) => data_im_in(505),
            data_re_out(0) => first_stage_re_out(25),
            data_re_out(1) => first_stage_re_out(57),
            data_re_out(2) => first_stage_re_out(89),
            data_re_out(3) => first_stage_re_out(121),
            data_re_out(4) => first_stage_re_out(153),
            data_re_out(5) => first_stage_re_out(185),
            data_re_out(6) => first_stage_re_out(217),
            data_re_out(7) => first_stage_re_out(249),
            data_re_out(8) => first_stage_re_out(281),
            data_re_out(9) => first_stage_re_out(313),
            data_re_out(10) => first_stage_re_out(345),
            data_re_out(11) => first_stage_re_out(377),
            data_re_out(12) => first_stage_re_out(409),
            data_re_out(13) => first_stage_re_out(441),
            data_re_out(14) => first_stage_re_out(473),
            data_re_out(15) => first_stage_re_out(505),
            data_im_out(0) => first_stage_im_out(25),
            data_im_out(1) => first_stage_im_out(57),
            data_im_out(2) => first_stage_im_out(89),
            data_im_out(3) => first_stage_im_out(121),
            data_im_out(4) => first_stage_im_out(153),
            data_im_out(5) => first_stage_im_out(185),
            data_im_out(6) => first_stage_im_out(217),
            data_im_out(7) => first_stage_im_out(249),
            data_im_out(8) => first_stage_im_out(281),
            data_im_out(9) => first_stage_im_out(313),
            data_im_out(10) => first_stage_im_out(345),
            data_im_out(11) => first_stage_im_out(377),
            data_im_out(12) => first_stage_im_out(409),
            data_im_out(13) => first_stage_im_out(441),
            data_im_out(14) => first_stage_im_out(473),
            data_im_out(15) => first_stage_im_out(505)
        );

    ULFFT_PT16_26 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(26),
            data_re_in(1) => data_re_in(58),
            data_re_in(2) => data_re_in(90),
            data_re_in(3) => data_re_in(122),
            data_re_in(4) => data_re_in(154),
            data_re_in(5) => data_re_in(186),
            data_re_in(6) => data_re_in(218),
            data_re_in(7) => data_re_in(250),
            data_re_in(8) => data_re_in(282),
            data_re_in(9) => data_re_in(314),
            data_re_in(10) => data_re_in(346),
            data_re_in(11) => data_re_in(378),
            data_re_in(12) => data_re_in(410),
            data_re_in(13) => data_re_in(442),
            data_re_in(14) => data_re_in(474),
            data_re_in(15) => data_re_in(506),
            data_im_in(0) => data_im_in(26),
            data_im_in(1) => data_im_in(58),
            data_im_in(2) => data_im_in(90),
            data_im_in(3) => data_im_in(122),
            data_im_in(4) => data_im_in(154),
            data_im_in(5) => data_im_in(186),
            data_im_in(6) => data_im_in(218),
            data_im_in(7) => data_im_in(250),
            data_im_in(8) => data_im_in(282),
            data_im_in(9) => data_im_in(314),
            data_im_in(10) => data_im_in(346),
            data_im_in(11) => data_im_in(378),
            data_im_in(12) => data_im_in(410),
            data_im_in(13) => data_im_in(442),
            data_im_in(14) => data_im_in(474),
            data_im_in(15) => data_im_in(506),
            data_re_out(0) => first_stage_re_out(26),
            data_re_out(1) => first_stage_re_out(58),
            data_re_out(2) => first_stage_re_out(90),
            data_re_out(3) => first_stage_re_out(122),
            data_re_out(4) => first_stage_re_out(154),
            data_re_out(5) => first_stage_re_out(186),
            data_re_out(6) => first_stage_re_out(218),
            data_re_out(7) => first_stage_re_out(250),
            data_re_out(8) => first_stage_re_out(282),
            data_re_out(9) => first_stage_re_out(314),
            data_re_out(10) => first_stage_re_out(346),
            data_re_out(11) => first_stage_re_out(378),
            data_re_out(12) => first_stage_re_out(410),
            data_re_out(13) => first_stage_re_out(442),
            data_re_out(14) => first_stage_re_out(474),
            data_re_out(15) => first_stage_re_out(506),
            data_im_out(0) => first_stage_im_out(26),
            data_im_out(1) => first_stage_im_out(58),
            data_im_out(2) => first_stage_im_out(90),
            data_im_out(3) => first_stage_im_out(122),
            data_im_out(4) => first_stage_im_out(154),
            data_im_out(5) => first_stage_im_out(186),
            data_im_out(6) => first_stage_im_out(218),
            data_im_out(7) => first_stage_im_out(250),
            data_im_out(8) => first_stage_im_out(282),
            data_im_out(9) => first_stage_im_out(314),
            data_im_out(10) => first_stage_im_out(346),
            data_im_out(11) => first_stage_im_out(378),
            data_im_out(12) => first_stage_im_out(410),
            data_im_out(13) => first_stage_im_out(442),
            data_im_out(14) => first_stage_im_out(474),
            data_im_out(15) => first_stage_im_out(506)
        );

    ULFFT_PT16_27 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(27),
            data_re_in(1) => data_re_in(59),
            data_re_in(2) => data_re_in(91),
            data_re_in(3) => data_re_in(123),
            data_re_in(4) => data_re_in(155),
            data_re_in(5) => data_re_in(187),
            data_re_in(6) => data_re_in(219),
            data_re_in(7) => data_re_in(251),
            data_re_in(8) => data_re_in(283),
            data_re_in(9) => data_re_in(315),
            data_re_in(10) => data_re_in(347),
            data_re_in(11) => data_re_in(379),
            data_re_in(12) => data_re_in(411),
            data_re_in(13) => data_re_in(443),
            data_re_in(14) => data_re_in(475),
            data_re_in(15) => data_re_in(507),
            data_im_in(0) => data_im_in(27),
            data_im_in(1) => data_im_in(59),
            data_im_in(2) => data_im_in(91),
            data_im_in(3) => data_im_in(123),
            data_im_in(4) => data_im_in(155),
            data_im_in(5) => data_im_in(187),
            data_im_in(6) => data_im_in(219),
            data_im_in(7) => data_im_in(251),
            data_im_in(8) => data_im_in(283),
            data_im_in(9) => data_im_in(315),
            data_im_in(10) => data_im_in(347),
            data_im_in(11) => data_im_in(379),
            data_im_in(12) => data_im_in(411),
            data_im_in(13) => data_im_in(443),
            data_im_in(14) => data_im_in(475),
            data_im_in(15) => data_im_in(507),
            data_re_out(0) => first_stage_re_out(27),
            data_re_out(1) => first_stage_re_out(59),
            data_re_out(2) => first_stage_re_out(91),
            data_re_out(3) => first_stage_re_out(123),
            data_re_out(4) => first_stage_re_out(155),
            data_re_out(5) => first_stage_re_out(187),
            data_re_out(6) => first_stage_re_out(219),
            data_re_out(7) => first_stage_re_out(251),
            data_re_out(8) => first_stage_re_out(283),
            data_re_out(9) => first_stage_re_out(315),
            data_re_out(10) => first_stage_re_out(347),
            data_re_out(11) => first_stage_re_out(379),
            data_re_out(12) => first_stage_re_out(411),
            data_re_out(13) => first_stage_re_out(443),
            data_re_out(14) => first_stage_re_out(475),
            data_re_out(15) => first_stage_re_out(507),
            data_im_out(0) => first_stage_im_out(27),
            data_im_out(1) => first_stage_im_out(59),
            data_im_out(2) => first_stage_im_out(91),
            data_im_out(3) => first_stage_im_out(123),
            data_im_out(4) => first_stage_im_out(155),
            data_im_out(5) => first_stage_im_out(187),
            data_im_out(6) => first_stage_im_out(219),
            data_im_out(7) => first_stage_im_out(251),
            data_im_out(8) => first_stage_im_out(283),
            data_im_out(9) => first_stage_im_out(315),
            data_im_out(10) => first_stage_im_out(347),
            data_im_out(11) => first_stage_im_out(379),
            data_im_out(12) => first_stage_im_out(411),
            data_im_out(13) => first_stage_im_out(443),
            data_im_out(14) => first_stage_im_out(475),
            data_im_out(15) => first_stage_im_out(507)
        );

    ULFFT_PT16_28 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(28),
            data_re_in(1) => data_re_in(60),
            data_re_in(2) => data_re_in(92),
            data_re_in(3) => data_re_in(124),
            data_re_in(4) => data_re_in(156),
            data_re_in(5) => data_re_in(188),
            data_re_in(6) => data_re_in(220),
            data_re_in(7) => data_re_in(252),
            data_re_in(8) => data_re_in(284),
            data_re_in(9) => data_re_in(316),
            data_re_in(10) => data_re_in(348),
            data_re_in(11) => data_re_in(380),
            data_re_in(12) => data_re_in(412),
            data_re_in(13) => data_re_in(444),
            data_re_in(14) => data_re_in(476),
            data_re_in(15) => data_re_in(508),
            data_im_in(0) => data_im_in(28),
            data_im_in(1) => data_im_in(60),
            data_im_in(2) => data_im_in(92),
            data_im_in(3) => data_im_in(124),
            data_im_in(4) => data_im_in(156),
            data_im_in(5) => data_im_in(188),
            data_im_in(6) => data_im_in(220),
            data_im_in(7) => data_im_in(252),
            data_im_in(8) => data_im_in(284),
            data_im_in(9) => data_im_in(316),
            data_im_in(10) => data_im_in(348),
            data_im_in(11) => data_im_in(380),
            data_im_in(12) => data_im_in(412),
            data_im_in(13) => data_im_in(444),
            data_im_in(14) => data_im_in(476),
            data_im_in(15) => data_im_in(508),
            data_re_out(0) => first_stage_re_out(28),
            data_re_out(1) => first_stage_re_out(60),
            data_re_out(2) => first_stage_re_out(92),
            data_re_out(3) => first_stage_re_out(124),
            data_re_out(4) => first_stage_re_out(156),
            data_re_out(5) => first_stage_re_out(188),
            data_re_out(6) => first_stage_re_out(220),
            data_re_out(7) => first_stage_re_out(252),
            data_re_out(8) => first_stage_re_out(284),
            data_re_out(9) => first_stage_re_out(316),
            data_re_out(10) => first_stage_re_out(348),
            data_re_out(11) => first_stage_re_out(380),
            data_re_out(12) => first_stage_re_out(412),
            data_re_out(13) => first_stage_re_out(444),
            data_re_out(14) => first_stage_re_out(476),
            data_re_out(15) => first_stage_re_out(508),
            data_im_out(0) => first_stage_im_out(28),
            data_im_out(1) => first_stage_im_out(60),
            data_im_out(2) => first_stage_im_out(92),
            data_im_out(3) => first_stage_im_out(124),
            data_im_out(4) => first_stage_im_out(156),
            data_im_out(5) => first_stage_im_out(188),
            data_im_out(6) => first_stage_im_out(220),
            data_im_out(7) => first_stage_im_out(252),
            data_im_out(8) => first_stage_im_out(284),
            data_im_out(9) => first_stage_im_out(316),
            data_im_out(10) => first_stage_im_out(348),
            data_im_out(11) => first_stage_im_out(380),
            data_im_out(12) => first_stage_im_out(412),
            data_im_out(13) => first_stage_im_out(444),
            data_im_out(14) => first_stage_im_out(476),
            data_im_out(15) => first_stage_im_out(508)
        );

    ULFFT_PT16_29 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(29),
            data_re_in(1) => data_re_in(61),
            data_re_in(2) => data_re_in(93),
            data_re_in(3) => data_re_in(125),
            data_re_in(4) => data_re_in(157),
            data_re_in(5) => data_re_in(189),
            data_re_in(6) => data_re_in(221),
            data_re_in(7) => data_re_in(253),
            data_re_in(8) => data_re_in(285),
            data_re_in(9) => data_re_in(317),
            data_re_in(10) => data_re_in(349),
            data_re_in(11) => data_re_in(381),
            data_re_in(12) => data_re_in(413),
            data_re_in(13) => data_re_in(445),
            data_re_in(14) => data_re_in(477),
            data_re_in(15) => data_re_in(509),
            data_im_in(0) => data_im_in(29),
            data_im_in(1) => data_im_in(61),
            data_im_in(2) => data_im_in(93),
            data_im_in(3) => data_im_in(125),
            data_im_in(4) => data_im_in(157),
            data_im_in(5) => data_im_in(189),
            data_im_in(6) => data_im_in(221),
            data_im_in(7) => data_im_in(253),
            data_im_in(8) => data_im_in(285),
            data_im_in(9) => data_im_in(317),
            data_im_in(10) => data_im_in(349),
            data_im_in(11) => data_im_in(381),
            data_im_in(12) => data_im_in(413),
            data_im_in(13) => data_im_in(445),
            data_im_in(14) => data_im_in(477),
            data_im_in(15) => data_im_in(509),
            data_re_out(0) => first_stage_re_out(29),
            data_re_out(1) => first_stage_re_out(61),
            data_re_out(2) => first_stage_re_out(93),
            data_re_out(3) => first_stage_re_out(125),
            data_re_out(4) => first_stage_re_out(157),
            data_re_out(5) => first_stage_re_out(189),
            data_re_out(6) => first_stage_re_out(221),
            data_re_out(7) => first_stage_re_out(253),
            data_re_out(8) => first_stage_re_out(285),
            data_re_out(9) => first_stage_re_out(317),
            data_re_out(10) => first_stage_re_out(349),
            data_re_out(11) => first_stage_re_out(381),
            data_re_out(12) => first_stage_re_out(413),
            data_re_out(13) => first_stage_re_out(445),
            data_re_out(14) => first_stage_re_out(477),
            data_re_out(15) => first_stage_re_out(509),
            data_im_out(0) => first_stage_im_out(29),
            data_im_out(1) => first_stage_im_out(61),
            data_im_out(2) => first_stage_im_out(93),
            data_im_out(3) => first_stage_im_out(125),
            data_im_out(4) => first_stage_im_out(157),
            data_im_out(5) => first_stage_im_out(189),
            data_im_out(6) => first_stage_im_out(221),
            data_im_out(7) => first_stage_im_out(253),
            data_im_out(8) => first_stage_im_out(285),
            data_im_out(9) => first_stage_im_out(317),
            data_im_out(10) => first_stage_im_out(349),
            data_im_out(11) => first_stage_im_out(381),
            data_im_out(12) => first_stage_im_out(413),
            data_im_out(13) => first_stage_im_out(445),
            data_im_out(14) => first_stage_im_out(477),
            data_im_out(15) => first_stage_im_out(509)
        );

    ULFFT_PT16_30 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(30),
            data_re_in(1) => data_re_in(62),
            data_re_in(2) => data_re_in(94),
            data_re_in(3) => data_re_in(126),
            data_re_in(4) => data_re_in(158),
            data_re_in(5) => data_re_in(190),
            data_re_in(6) => data_re_in(222),
            data_re_in(7) => data_re_in(254),
            data_re_in(8) => data_re_in(286),
            data_re_in(9) => data_re_in(318),
            data_re_in(10) => data_re_in(350),
            data_re_in(11) => data_re_in(382),
            data_re_in(12) => data_re_in(414),
            data_re_in(13) => data_re_in(446),
            data_re_in(14) => data_re_in(478),
            data_re_in(15) => data_re_in(510),
            data_im_in(0) => data_im_in(30),
            data_im_in(1) => data_im_in(62),
            data_im_in(2) => data_im_in(94),
            data_im_in(3) => data_im_in(126),
            data_im_in(4) => data_im_in(158),
            data_im_in(5) => data_im_in(190),
            data_im_in(6) => data_im_in(222),
            data_im_in(7) => data_im_in(254),
            data_im_in(8) => data_im_in(286),
            data_im_in(9) => data_im_in(318),
            data_im_in(10) => data_im_in(350),
            data_im_in(11) => data_im_in(382),
            data_im_in(12) => data_im_in(414),
            data_im_in(13) => data_im_in(446),
            data_im_in(14) => data_im_in(478),
            data_im_in(15) => data_im_in(510),
            data_re_out(0) => first_stage_re_out(30),
            data_re_out(1) => first_stage_re_out(62),
            data_re_out(2) => first_stage_re_out(94),
            data_re_out(3) => first_stage_re_out(126),
            data_re_out(4) => first_stage_re_out(158),
            data_re_out(5) => first_stage_re_out(190),
            data_re_out(6) => first_stage_re_out(222),
            data_re_out(7) => first_stage_re_out(254),
            data_re_out(8) => first_stage_re_out(286),
            data_re_out(9) => first_stage_re_out(318),
            data_re_out(10) => first_stage_re_out(350),
            data_re_out(11) => first_stage_re_out(382),
            data_re_out(12) => first_stage_re_out(414),
            data_re_out(13) => first_stage_re_out(446),
            data_re_out(14) => first_stage_re_out(478),
            data_re_out(15) => first_stage_re_out(510),
            data_im_out(0) => first_stage_im_out(30),
            data_im_out(1) => first_stage_im_out(62),
            data_im_out(2) => first_stage_im_out(94),
            data_im_out(3) => first_stage_im_out(126),
            data_im_out(4) => first_stage_im_out(158),
            data_im_out(5) => first_stage_im_out(190),
            data_im_out(6) => first_stage_im_out(222),
            data_im_out(7) => first_stage_im_out(254),
            data_im_out(8) => first_stage_im_out(286),
            data_im_out(9) => first_stage_im_out(318),
            data_im_out(10) => first_stage_im_out(350),
            data_im_out(11) => first_stage_im_out(382),
            data_im_out(12) => first_stage_im_out(414),
            data_im_out(13) => first_stage_im_out(446),
            data_im_out(14) => first_stage_im_out(478),
            data_im_out(15) => first_stage_im_out(510)
        );

    ULFFT_PT16_31 : fft_pt16
    generic map(
        ctrl_start => ctrl_start
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(8 DOWNTO 5),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => data_re_in(31),
            data_re_in(1) => data_re_in(63),
            data_re_in(2) => data_re_in(95),
            data_re_in(3) => data_re_in(127),
            data_re_in(4) => data_re_in(159),
            data_re_in(5) => data_re_in(191),
            data_re_in(6) => data_re_in(223),
            data_re_in(7) => data_re_in(255),
            data_re_in(8) => data_re_in(287),
            data_re_in(9) => data_re_in(319),
            data_re_in(10) => data_re_in(351),
            data_re_in(11) => data_re_in(383),
            data_re_in(12) => data_re_in(415),
            data_re_in(13) => data_re_in(447),
            data_re_in(14) => data_re_in(479),
            data_re_in(15) => data_re_in(511),
            data_im_in(0) => data_im_in(31),
            data_im_in(1) => data_im_in(63),
            data_im_in(2) => data_im_in(95),
            data_im_in(3) => data_im_in(127),
            data_im_in(4) => data_im_in(159),
            data_im_in(5) => data_im_in(191),
            data_im_in(6) => data_im_in(223),
            data_im_in(7) => data_im_in(255),
            data_im_in(8) => data_im_in(287),
            data_im_in(9) => data_im_in(319),
            data_im_in(10) => data_im_in(351),
            data_im_in(11) => data_im_in(383),
            data_im_in(12) => data_im_in(415),
            data_im_in(13) => data_im_in(447),
            data_im_in(14) => data_im_in(479),
            data_im_in(15) => data_im_in(511),
            data_re_out(0) => first_stage_re_out(31),
            data_re_out(1) => first_stage_re_out(63),
            data_re_out(2) => first_stage_re_out(95),
            data_re_out(3) => first_stage_re_out(127),
            data_re_out(4) => first_stage_re_out(159),
            data_re_out(5) => first_stage_re_out(191),
            data_re_out(6) => first_stage_re_out(223),
            data_re_out(7) => first_stage_re_out(255),
            data_re_out(8) => first_stage_re_out(287),
            data_re_out(9) => first_stage_re_out(319),
            data_re_out(10) => first_stage_re_out(351),
            data_re_out(11) => first_stage_re_out(383),
            data_re_out(12) => first_stage_re_out(415),
            data_re_out(13) => first_stage_re_out(447),
            data_re_out(14) => first_stage_re_out(479),
            data_re_out(15) => first_stage_re_out(511),
            data_im_out(0) => first_stage_im_out(31),
            data_im_out(1) => first_stage_im_out(63),
            data_im_out(2) => first_stage_im_out(95),
            data_im_out(3) => first_stage_im_out(127),
            data_im_out(4) => first_stage_im_out(159),
            data_im_out(5) => first_stage_im_out(191),
            data_im_out(6) => first_stage_im_out(223),
            data_im_out(7) => first_stage_im_out(255),
            data_im_out(8) => first_stage_im_out(287),
            data_im_out(9) => first_stage_im_out(319),
            data_im_out(10) => first_stage_im_out(351),
            data_im_out(11) => first_stage_im_out(383),
            data_im_out(12) => first_stage_im_out(415),
            data_im_out(13) => first_stage_im_out(447),
            data_im_out(14) => first_stage_im_out(479),
            data_im_out(15) => first_stage_im_out(511)
        );


    --- right-hand-side processors
    URFFT_PT32_0 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(0),
            data_re_in(1) => mul_re_out(1),
            data_re_in(2) => mul_re_out(2),
            data_re_in(3) => mul_re_out(3),
            data_re_in(4) => mul_re_out(4),
            data_re_in(5) => mul_re_out(5),
            data_re_in(6) => mul_re_out(6),
            data_re_in(7) => mul_re_out(7),
            data_re_in(8) => mul_re_out(8),
            data_re_in(9) => mul_re_out(9),
            data_re_in(10) => mul_re_out(10),
            data_re_in(11) => mul_re_out(11),
            data_re_in(12) => mul_re_out(12),
            data_re_in(13) => mul_re_out(13),
            data_re_in(14) => mul_re_out(14),
            data_re_in(15) => mul_re_out(15),
            data_re_in(16) => mul_re_out(16),
            data_re_in(17) => mul_re_out(17),
            data_re_in(18) => mul_re_out(18),
            data_re_in(19) => mul_re_out(19),
            data_re_in(20) => mul_re_out(20),
            data_re_in(21) => mul_re_out(21),
            data_re_in(22) => mul_re_out(22),
            data_re_in(23) => mul_re_out(23),
            data_re_in(24) => mul_re_out(24),
            data_re_in(25) => mul_re_out(25),
            data_re_in(26) => mul_re_out(26),
            data_re_in(27) => mul_re_out(27),
            data_re_in(28) => mul_re_out(28),
            data_re_in(29) => mul_re_out(29),
            data_re_in(30) => mul_re_out(30),
            data_re_in(31) => mul_re_out(31),
            data_im_in(0) => mul_im_out(0),
            data_im_in(1) => mul_im_out(1),
            data_im_in(2) => mul_im_out(2),
            data_im_in(3) => mul_im_out(3),
            data_im_in(4) => mul_im_out(4),
            data_im_in(5) => mul_im_out(5),
            data_im_in(6) => mul_im_out(6),
            data_im_in(7) => mul_im_out(7),
            data_im_in(8) => mul_im_out(8),
            data_im_in(9) => mul_im_out(9),
            data_im_in(10) => mul_im_out(10),
            data_im_in(11) => mul_im_out(11),
            data_im_in(12) => mul_im_out(12),
            data_im_in(13) => mul_im_out(13),
            data_im_in(14) => mul_im_out(14),
            data_im_in(15) => mul_im_out(15),
            data_im_in(16) => mul_im_out(16),
            data_im_in(17) => mul_im_out(17),
            data_im_in(18) => mul_im_out(18),
            data_im_in(19) => mul_im_out(19),
            data_im_in(20) => mul_im_out(20),
            data_im_in(21) => mul_im_out(21),
            data_im_in(22) => mul_im_out(22),
            data_im_in(23) => mul_im_out(23),
            data_im_in(24) => mul_im_out(24),
            data_im_in(25) => mul_im_out(25),
            data_im_in(26) => mul_im_out(26),
            data_im_in(27) => mul_im_out(27),
            data_im_in(28) => mul_im_out(28),
            data_im_in(29) => mul_im_out(29),
            data_im_in(30) => mul_im_out(30),
            data_im_in(31) => mul_im_out(31),
            data_re_out(0) => data_re_out(0),
            data_re_out(1) => data_re_out(16),
            data_re_out(2) => data_re_out(32),
            data_re_out(3) => data_re_out(48),
            data_re_out(4) => data_re_out(64),
            data_re_out(5) => data_re_out(80),
            data_re_out(6) => data_re_out(96),
            data_re_out(7) => data_re_out(112),
            data_re_out(8) => data_re_out(128),
            data_re_out(9) => data_re_out(144),
            data_re_out(10) => data_re_out(160),
            data_re_out(11) => data_re_out(176),
            data_re_out(12) => data_re_out(192),
            data_re_out(13) => data_re_out(208),
            data_re_out(14) => data_re_out(224),
            data_re_out(15) => data_re_out(240),
            data_re_out(16) => data_re_out(256),
            data_re_out(17) => data_re_out(272),
            data_re_out(18) => data_re_out(288),
            data_re_out(19) => data_re_out(304),
            data_re_out(20) => data_re_out(320),
            data_re_out(21) => data_re_out(336),
            data_re_out(22) => data_re_out(352),
            data_re_out(23) => data_re_out(368),
            data_re_out(24) => data_re_out(384),
            data_re_out(25) => data_re_out(400),
            data_re_out(26) => data_re_out(416),
            data_re_out(27) => data_re_out(432),
            data_re_out(28) => data_re_out(448),
            data_re_out(29) => data_re_out(464),
            data_re_out(30) => data_re_out(480),
            data_re_out(31) => data_re_out(496),
            data_im_out(0) => data_im_out(0),
            data_im_out(1) => data_im_out(16),
            data_im_out(2) => data_im_out(32),
            data_im_out(3) => data_im_out(48),
            data_im_out(4) => data_im_out(64),
            data_im_out(5) => data_im_out(80),
            data_im_out(6) => data_im_out(96),
            data_im_out(7) => data_im_out(112),
            data_im_out(8) => data_im_out(128),
            data_im_out(9) => data_im_out(144),
            data_im_out(10) => data_im_out(160),
            data_im_out(11) => data_im_out(176),
            data_im_out(12) => data_im_out(192),
            data_im_out(13) => data_im_out(208),
            data_im_out(14) => data_im_out(224),
            data_im_out(15) => data_im_out(240),
            data_im_out(16) => data_im_out(256),
            data_im_out(17) => data_im_out(272),
            data_im_out(18) => data_im_out(288),
            data_im_out(19) => data_im_out(304),
            data_im_out(20) => data_im_out(320),
            data_im_out(21) => data_im_out(336),
            data_im_out(22) => data_im_out(352),
            data_im_out(23) => data_im_out(368),
            data_im_out(24) => data_im_out(384),
            data_im_out(25) => data_im_out(400),
            data_im_out(26) => data_im_out(416),
            data_im_out(27) => data_im_out(432),
            data_im_out(28) => data_im_out(448),
            data_im_out(29) => data_im_out(464),
            data_im_out(30) => data_im_out(480),
            data_im_out(31) => data_im_out(496)
        );           

    URFFT_PT32_1 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(32),
            data_re_in(1) => mul_re_out(33),
            data_re_in(2) => mul_re_out(34),
            data_re_in(3) => mul_re_out(35),
            data_re_in(4) => mul_re_out(36),
            data_re_in(5) => mul_re_out(37),
            data_re_in(6) => mul_re_out(38),
            data_re_in(7) => mul_re_out(39),
            data_re_in(8) => mul_re_out(40),
            data_re_in(9) => mul_re_out(41),
            data_re_in(10) => mul_re_out(42),
            data_re_in(11) => mul_re_out(43),
            data_re_in(12) => mul_re_out(44),
            data_re_in(13) => mul_re_out(45),
            data_re_in(14) => mul_re_out(46),
            data_re_in(15) => mul_re_out(47),
            data_re_in(16) => mul_re_out(48),
            data_re_in(17) => mul_re_out(49),
            data_re_in(18) => mul_re_out(50),
            data_re_in(19) => mul_re_out(51),
            data_re_in(20) => mul_re_out(52),
            data_re_in(21) => mul_re_out(53),
            data_re_in(22) => mul_re_out(54),
            data_re_in(23) => mul_re_out(55),
            data_re_in(24) => mul_re_out(56),
            data_re_in(25) => mul_re_out(57),
            data_re_in(26) => mul_re_out(58),
            data_re_in(27) => mul_re_out(59),
            data_re_in(28) => mul_re_out(60),
            data_re_in(29) => mul_re_out(61),
            data_re_in(30) => mul_re_out(62),
            data_re_in(31) => mul_re_out(63),
            data_im_in(0) => mul_im_out(32),
            data_im_in(1) => mul_im_out(33),
            data_im_in(2) => mul_im_out(34),
            data_im_in(3) => mul_im_out(35),
            data_im_in(4) => mul_im_out(36),
            data_im_in(5) => mul_im_out(37),
            data_im_in(6) => mul_im_out(38),
            data_im_in(7) => mul_im_out(39),
            data_im_in(8) => mul_im_out(40),
            data_im_in(9) => mul_im_out(41),
            data_im_in(10) => mul_im_out(42),
            data_im_in(11) => mul_im_out(43),
            data_im_in(12) => mul_im_out(44),
            data_im_in(13) => mul_im_out(45),
            data_im_in(14) => mul_im_out(46),
            data_im_in(15) => mul_im_out(47),
            data_im_in(16) => mul_im_out(48),
            data_im_in(17) => mul_im_out(49),
            data_im_in(18) => mul_im_out(50),
            data_im_in(19) => mul_im_out(51),
            data_im_in(20) => mul_im_out(52),
            data_im_in(21) => mul_im_out(53),
            data_im_in(22) => mul_im_out(54),
            data_im_in(23) => mul_im_out(55),
            data_im_in(24) => mul_im_out(56),
            data_im_in(25) => mul_im_out(57),
            data_im_in(26) => mul_im_out(58),
            data_im_in(27) => mul_im_out(59),
            data_im_in(28) => mul_im_out(60),
            data_im_in(29) => mul_im_out(61),
            data_im_in(30) => mul_im_out(62),
            data_im_in(31) => mul_im_out(63),
            data_re_out(0) => data_re_out(1),
            data_re_out(1) => data_re_out(17),
            data_re_out(2) => data_re_out(33),
            data_re_out(3) => data_re_out(49),
            data_re_out(4) => data_re_out(65),
            data_re_out(5) => data_re_out(81),
            data_re_out(6) => data_re_out(97),
            data_re_out(7) => data_re_out(113),
            data_re_out(8) => data_re_out(129),
            data_re_out(9) => data_re_out(145),
            data_re_out(10) => data_re_out(161),
            data_re_out(11) => data_re_out(177),
            data_re_out(12) => data_re_out(193),
            data_re_out(13) => data_re_out(209),
            data_re_out(14) => data_re_out(225),
            data_re_out(15) => data_re_out(241),
            data_re_out(16) => data_re_out(257),
            data_re_out(17) => data_re_out(273),
            data_re_out(18) => data_re_out(289),
            data_re_out(19) => data_re_out(305),
            data_re_out(20) => data_re_out(321),
            data_re_out(21) => data_re_out(337),
            data_re_out(22) => data_re_out(353),
            data_re_out(23) => data_re_out(369),
            data_re_out(24) => data_re_out(385),
            data_re_out(25) => data_re_out(401),
            data_re_out(26) => data_re_out(417),
            data_re_out(27) => data_re_out(433),
            data_re_out(28) => data_re_out(449),
            data_re_out(29) => data_re_out(465),
            data_re_out(30) => data_re_out(481),
            data_re_out(31) => data_re_out(497),
            data_im_out(0) => data_im_out(1),
            data_im_out(1) => data_im_out(17),
            data_im_out(2) => data_im_out(33),
            data_im_out(3) => data_im_out(49),
            data_im_out(4) => data_im_out(65),
            data_im_out(5) => data_im_out(81),
            data_im_out(6) => data_im_out(97),
            data_im_out(7) => data_im_out(113),
            data_im_out(8) => data_im_out(129),
            data_im_out(9) => data_im_out(145),
            data_im_out(10) => data_im_out(161),
            data_im_out(11) => data_im_out(177),
            data_im_out(12) => data_im_out(193),
            data_im_out(13) => data_im_out(209),
            data_im_out(14) => data_im_out(225),
            data_im_out(15) => data_im_out(241),
            data_im_out(16) => data_im_out(257),
            data_im_out(17) => data_im_out(273),
            data_im_out(18) => data_im_out(289),
            data_im_out(19) => data_im_out(305),
            data_im_out(20) => data_im_out(321),
            data_im_out(21) => data_im_out(337),
            data_im_out(22) => data_im_out(353),
            data_im_out(23) => data_im_out(369),
            data_im_out(24) => data_im_out(385),
            data_im_out(25) => data_im_out(401),
            data_im_out(26) => data_im_out(417),
            data_im_out(27) => data_im_out(433),
            data_im_out(28) => data_im_out(449),
            data_im_out(29) => data_im_out(465),
            data_im_out(30) => data_im_out(481),
            data_im_out(31) => data_im_out(497)
        );           

    URFFT_PT32_2 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(64),
            data_re_in(1) => mul_re_out(65),
            data_re_in(2) => mul_re_out(66),
            data_re_in(3) => mul_re_out(67),
            data_re_in(4) => mul_re_out(68),
            data_re_in(5) => mul_re_out(69),
            data_re_in(6) => mul_re_out(70),
            data_re_in(7) => mul_re_out(71),
            data_re_in(8) => mul_re_out(72),
            data_re_in(9) => mul_re_out(73),
            data_re_in(10) => mul_re_out(74),
            data_re_in(11) => mul_re_out(75),
            data_re_in(12) => mul_re_out(76),
            data_re_in(13) => mul_re_out(77),
            data_re_in(14) => mul_re_out(78),
            data_re_in(15) => mul_re_out(79),
            data_re_in(16) => mul_re_out(80),
            data_re_in(17) => mul_re_out(81),
            data_re_in(18) => mul_re_out(82),
            data_re_in(19) => mul_re_out(83),
            data_re_in(20) => mul_re_out(84),
            data_re_in(21) => mul_re_out(85),
            data_re_in(22) => mul_re_out(86),
            data_re_in(23) => mul_re_out(87),
            data_re_in(24) => mul_re_out(88),
            data_re_in(25) => mul_re_out(89),
            data_re_in(26) => mul_re_out(90),
            data_re_in(27) => mul_re_out(91),
            data_re_in(28) => mul_re_out(92),
            data_re_in(29) => mul_re_out(93),
            data_re_in(30) => mul_re_out(94),
            data_re_in(31) => mul_re_out(95),
            data_im_in(0) => mul_im_out(64),
            data_im_in(1) => mul_im_out(65),
            data_im_in(2) => mul_im_out(66),
            data_im_in(3) => mul_im_out(67),
            data_im_in(4) => mul_im_out(68),
            data_im_in(5) => mul_im_out(69),
            data_im_in(6) => mul_im_out(70),
            data_im_in(7) => mul_im_out(71),
            data_im_in(8) => mul_im_out(72),
            data_im_in(9) => mul_im_out(73),
            data_im_in(10) => mul_im_out(74),
            data_im_in(11) => mul_im_out(75),
            data_im_in(12) => mul_im_out(76),
            data_im_in(13) => mul_im_out(77),
            data_im_in(14) => mul_im_out(78),
            data_im_in(15) => mul_im_out(79),
            data_im_in(16) => mul_im_out(80),
            data_im_in(17) => mul_im_out(81),
            data_im_in(18) => mul_im_out(82),
            data_im_in(19) => mul_im_out(83),
            data_im_in(20) => mul_im_out(84),
            data_im_in(21) => mul_im_out(85),
            data_im_in(22) => mul_im_out(86),
            data_im_in(23) => mul_im_out(87),
            data_im_in(24) => mul_im_out(88),
            data_im_in(25) => mul_im_out(89),
            data_im_in(26) => mul_im_out(90),
            data_im_in(27) => mul_im_out(91),
            data_im_in(28) => mul_im_out(92),
            data_im_in(29) => mul_im_out(93),
            data_im_in(30) => mul_im_out(94),
            data_im_in(31) => mul_im_out(95),
            data_re_out(0) => data_re_out(2),
            data_re_out(1) => data_re_out(18),
            data_re_out(2) => data_re_out(34),
            data_re_out(3) => data_re_out(50),
            data_re_out(4) => data_re_out(66),
            data_re_out(5) => data_re_out(82),
            data_re_out(6) => data_re_out(98),
            data_re_out(7) => data_re_out(114),
            data_re_out(8) => data_re_out(130),
            data_re_out(9) => data_re_out(146),
            data_re_out(10) => data_re_out(162),
            data_re_out(11) => data_re_out(178),
            data_re_out(12) => data_re_out(194),
            data_re_out(13) => data_re_out(210),
            data_re_out(14) => data_re_out(226),
            data_re_out(15) => data_re_out(242),
            data_re_out(16) => data_re_out(258),
            data_re_out(17) => data_re_out(274),
            data_re_out(18) => data_re_out(290),
            data_re_out(19) => data_re_out(306),
            data_re_out(20) => data_re_out(322),
            data_re_out(21) => data_re_out(338),
            data_re_out(22) => data_re_out(354),
            data_re_out(23) => data_re_out(370),
            data_re_out(24) => data_re_out(386),
            data_re_out(25) => data_re_out(402),
            data_re_out(26) => data_re_out(418),
            data_re_out(27) => data_re_out(434),
            data_re_out(28) => data_re_out(450),
            data_re_out(29) => data_re_out(466),
            data_re_out(30) => data_re_out(482),
            data_re_out(31) => data_re_out(498),
            data_im_out(0) => data_im_out(2),
            data_im_out(1) => data_im_out(18),
            data_im_out(2) => data_im_out(34),
            data_im_out(3) => data_im_out(50),
            data_im_out(4) => data_im_out(66),
            data_im_out(5) => data_im_out(82),
            data_im_out(6) => data_im_out(98),
            data_im_out(7) => data_im_out(114),
            data_im_out(8) => data_im_out(130),
            data_im_out(9) => data_im_out(146),
            data_im_out(10) => data_im_out(162),
            data_im_out(11) => data_im_out(178),
            data_im_out(12) => data_im_out(194),
            data_im_out(13) => data_im_out(210),
            data_im_out(14) => data_im_out(226),
            data_im_out(15) => data_im_out(242),
            data_im_out(16) => data_im_out(258),
            data_im_out(17) => data_im_out(274),
            data_im_out(18) => data_im_out(290),
            data_im_out(19) => data_im_out(306),
            data_im_out(20) => data_im_out(322),
            data_im_out(21) => data_im_out(338),
            data_im_out(22) => data_im_out(354),
            data_im_out(23) => data_im_out(370),
            data_im_out(24) => data_im_out(386),
            data_im_out(25) => data_im_out(402),
            data_im_out(26) => data_im_out(418),
            data_im_out(27) => data_im_out(434),
            data_im_out(28) => data_im_out(450),
            data_im_out(29) => data_im_out(466),
            data_im_out(30) => data_im_out(482),
            data_im_out(31) => data_im_out(498)
        );           

    URFFT_PT32_3 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(96),
            data_re_in(1) => mul_re_out(97),
            data_re_in(2) => mul_re_out(98),
            data_re_in(3) => mul_re_out(99),
            data_re_in(4) => mul_re_out(100),
            data_re_in(5) => mul_re_out(101),
            data_re_in(6) => mul_re_out(102),
            data_re_in(7) => mul_re_out(103),
            data_re_in(8) => mul_re_out(104),
            data_re_in(9) => mul_re_out(105),
            data_re_in(10) => mul_re_out(106),
            data_re_in(11) => mul_re_out(107),
            data_re_in(12) => mul_re_out(108),
            data_re_in(13) => mul_re_out(109),
            data_re_in(14) => mul_re_out(110),
            data_re_in(15) => mul_re_out(111),
            data_re_in(16) => mul_re_out(112),
            data_re_in(17) => mul_re_out(113),
            data_re_in(18) => mul_re_out(114),
            data_re_in(19) => mul_re_out(115),
            data_re_in(20) => mul_re_out(116),
            data_re_in(21) => mul_re_out(117),
            data_re_in(22) => mul_re_out(118),
            data_re_in(23) => mul_re_out(119),
            data_re_in(24) => mul_re_out(120),
            data_re_in(25) => mul_re_out(121),
            data_re_in(26) => mul_re_out(122),
            data_re_in(27) => mul_re_out(123),
            data_re_in(28) => mul_re_out(124),
            data_re_in(29) => mul_re_out(125),
            data_re_in(30) => mul_re_out(126),
            data_re_in(31) => mul_re_out(127),
            data_im_in(0) => mul_im_out(96),
            data_im_in(1) => mul_im_out(97),
            data_im_in(2) => mul_im_out(98),
            data_im_in(3) => mul_im_out(99),
            data_im_in(4) => mul_im_out(100),
            data_im_in(5) => mul_im_out(101),
            data_im_in(6) => mul_im_out(102),
            data_im_in(7) => mul_im_out(103),
            data_im_in(8) => mul_im_out(104),
            data_im_in(9) => mul_im_out(105),
            data_im_in(10) => mul_im_out(106),
            data_im_in(11) => mul_im_out(107),
            data_im_in(12) => mul_im_out(108),
            data_im_in(13) => mul_im_out(109),
            data_im_in(14) => mul_im_out(110),
            data_im_in(15) => mul_im_out(111),
            data_im_in(16) => mul_im_out(112),
            data_im_in(17) => mul_im_out(113),
            data_im_in(18) => mul_im_out(114),
            data_im_in(19) => mul_im_out(115),
            data_im_in(20) => mul_im_out(116),
            data_im_in(21) => mul_im_out(117),
            data_im_in(22) => mul_im_out(118),
            data_im_in(23) => mul_im_out(119),
            data_im_in(24) => mul_im_out(120),
            data_im_in(25) => mul_im_out(121),
            data_im_in(26) => mul_im_out(122),
            data_im_in(27) => mul_im_out(123),
            data_im_in(28) => mul_im_out(124),
            data_im_in(29) => mul_im_out(125),
            data_im_in(30) => mul_im_out(126),
            data_im_in(31) => mul_im_out(127),
            data_re_out(0) => data_re_out(3),
            data_re_out(1) => data_re_out(19),
            data_re_out(2) => data_re_out(35),
            data_re_out(3) => data_re_out(51),
            data_re_out(4) => data_re_out(67),
            data_re_out(5) => data_re_out(83),
            data_re_out(6) => data_re_out(99),
            data_re_out(7) => data_re_out(115),
            data_re_out(8) => data_re_out(131),
            data_re_out(9) => data_re_out(147),
            data_re_out(10) => data_re_out(163),
            data_re_out(11) => data_re_out(179),
            data_re_out(12) => data_re_out(195),
            data_re_out(13) => data_re_out(211),
            data_re_out(14) => data_re_out(227),
            data_re_out(15) => data_re_out(243),
            data_re_out(16) => data_re_out(259),
            data_re_out(17) => data_re_out(275),
            data_re_out(18) => data_re_out(291),
            data_re_out(19) => data_re_out(307),
            data_re_out(20) => data_re_out(323),
            data_re_out(21) => data_re_out(339),
            data_re_out(22) => data_re_out(355),
            data_re_out(23) => data_re_out(371),
            data_re_out(24) => data_re_out(387),
            data_re_out(25) => data_re_out(403),
            data_re_out(26) => data_re_out(419),
            data_re_out(27) => data_re_out(435),
            data_re_out(28) => data_re_out(451),
            data_re_out(29) => data_re_out(467),
            data_re_out(30) => data_re_out(483),
            data_re_out(31) => data_re_out(499),
            data_im_out(0) => data_im_out(3),
            data_im_out(1) => data_im_out(19),
            data_im_out(2) => data_im_out(35),
            data_im_out(3) => data_im_out(51),
            data_im_out(4) => data_im_out(67),
            data_im_out(5) => data_im_out(83),
            data_im_out(6) => data_im_out(99),
            data_im_out(7) => data_im_out(115),
            data_im_out(8) => data_im_out(131),
            data_im_out(9) => data_im_out(147),
            data_im_out(10) => data_im_out(163),
            data_im_out(11) => data_im_out(179),
            data_im_out(12) => data_im_out(195),
            data_im_out(13) => data_im_out(211),
            data_im_out(14) => data_im_out(227),
            data_im_out(15) => data_im_out(243),
            data_im_out(16) => data_im_out(259),
            data_im_out(17) => data_im_out(275),
            data_im_out(18) => data_im_out(291),
            data_im_out(19) => data_im_out(307),
            data_im_out(20) => data_im_out(323),
            data_im_out(21) => data_im_out(339),
            data_im_out(22) => data_im_out(355),
            data_im_out(23) => data_im_out(371),
            data_im_out(24) => data_im_out(387),
            data_im_out(25) => data_im_out(403),
            data_im_out(26) => data_im_out(419),
            data_im_out(27) => data_im_out(435),
            data_im_out(28) => data_im_out(451),
            data_im_out(29) => data_im_out(467),
            data_im_out(30) => data_im_out(483),
            data_im_out(31) => data_im_out(499)
        );           

    URFFT_PT32_4 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(128),
            data_re_in(1) => mul_re_out(129),
            data_re_in(2) => mul_re_out(130),
            data_re_in(3) => mul_re_out(131),
            data_re_in(4) => mul_re_out(132),
            data_re_in(5) => mul_re_out(133),
            data_re_in(6) => mul_re_out(134),
            data_re_in(7) => mul_re_out(135),
            data_re_in(8) => mul_re_out(136),
            data_re_in(9) => mul_re_out(137),
            data_re_in(10) => mul_re_out(138),
            data_re_in(11) => mul_re_out(139),
            data_re_in(12) => mul_re_out(140),
            data_re_in(13) => mul_re_out(141),
            data_re_in(14) => mul_re_out(142),
            data_re_in(15) => mul_re_out(143),
            data_re_in(16) => mul_re_out(144),
            data_re_in(17) => mul_re_out(145),
            data_re_in(18) => mul_re_out(146),
            data_re_in(19) => mul_re_out(147),
            data_re_in(20) => mul_re_out(148),
            data_re_in(21) => mul_re_out(149),
            data_re_in(22) => mul_re_out(150),
            data_re_in(23) => mul_re_out(151),
            data_re_in(24) => mul_re_out(152),
            data_re_in(25) => mul_re_out(153),
            data_re_in(26) => mul_re_out(154),
            data_re_in(27) => mul_re_out(155),
            data_re_in(28) => mul_re_out(156),
            data_re_in(29) => mul_re_out(157),
            data_re_in(30) => mul_re_out(158),
            data_re_in(31) => mul_re_out(159),
            data_im_in(0) => mul_im_out(128),
            data_im_in(1) => mul_im_out(129),
            data_im_in(2) => mul_im_out(130),
            data_im_in(3) => mul_im_out(131),
            data_im_in(4) => mul_im_out(132),
            data_im_in(5) => mul_im_out(133),
            data_im_in(6) => mul_im_out(134),
            data_im_in(7) => mul_im_out(135),
            data_im_in(8) => mul_im_out(136),
            data_im_in(9) => mul_im_out(137),
            data_im_in(10) => mul_im_out(138),
            data_im_in(11) => mul_im_out(139),
            data_im_in(12) => mul_im_out(140),
            data_im_in(13) => mul_im_out(141),
            data_im_in(14) => mul_im_out(142),
            data_im_in(15) => mul_im_out(143),
            data_im_in(16) => mul_im_out(144),
            data_im_in(17) => mul_im_out(145),
            data_im_in(18) => mul_im_out(146),
            data_im_in(19) => mul_im_out(147),
            data_im_in(20) => mul_im_out(148),
            data_im_in(21) => mul_im_out(149),
            data_im_in(22) => mul_im_out(150),
            data_im_in(23) => mul_im_out(151),
            data_im_in(24) => mul_im_out(152),
            data_im_in(25) => mul_im_out(153),
            data_im_in(26) => mul_im_out(154),
            data_im_in(27) => mul_im_out(155),
            data_im_in(28) => mul_im_out(156),
            data_im_in(29) => mul_im_out(157),
            data_im_in(30) => mul_im_out(158),
            data_im_in(31) => mul_im_out(159),
            data_re_out(0) => data_re_out(4),
            data_re_out(1) => data_re_out(20),
            data_re_out(2) => data_re_out(36),
            data_re_out(3) => data_re_out(52),
            data_re_out(4) => data_re_out(68),
            data_re_out(5) => data_re_out(84),
            data_re_out(6) => data_re_out(100),
            data_re_out(7) => data_re_out(116),
            data_re_out(8) => data_re_out(132),
            data_re_out(9) => data_re_out(148),
            data_re_out(10) => data_re_out(164),
            data_re_out(11) => data_re_out(180),
            data_re_out(12) => data_re_out(196),
            data_re_out(13) => data_re_out(212),
            data_re_out(14) => data_re_out(228),
            data_re_out(15) => data_re_out(244),
            data_re_out(16) => data_re_out(260),
            data_re_out(17) => data_re_out(276),
            data_re_out(18) => data_re_out(292),
            data_re_out(19) => data_re_out(308),
            data_re_out(20) => data_re_out(324),
            data_re_out(21) => data_re_out(340),
            data_re_out(22) => data_re_out(356),
            data_re_out(23) => data_re_out(372),
            data_re_out(24) => data_re_out(388),
            data_re_out(25) => data_re_out(404),
            data_re_out(26) => data_re_out(420),
            data_re_out(27) => data_re_out(436),
            data_re_out(28) => data_re_out(452),
            data_re_out(29) => data_re_out(468),
            data_re_out(30) => data_re_out(484),
            data_re_out(31) => data_re_out(500),
            data_im_out(0) => data_im_out(4),
            data_im_out(1) => data_im_out(20),
            data_im_out(2) => data_im_out(36),
            data_im_out(3) => data_im_out(52),
            data_im_out(4) => data_im_out(68),
            data_im_out(5) => data_im_out(84),
            data_im_out(6) => data_im_out(100),
            data_im_out(7) => data_im_out(116),
            data_im_out(8) => data_im_out(132),
            data_im_out(9) => data_im_out(148),
            data_im_out(10) => data_im_out(164),
            data_im_out(11) => data_im_out(180),
            data_im_out(12) => data_im_out(196),
            data_im_out(13) => data_im_out(212),
            data_im_out(14) => data_im_out(228),
            data_im_out(15) => data_im_out(244),
            data_im_out(16) => data_im_out(260),
            data_im_out(17) => data_im_out(276),
            data_im_out(18) => data_im_out(292),
            data_im_out(19) => data_im_out(308),
            data_im_out(20) => data_im_out(324),
            data_im_out(21) => data_im_out(340),
            data_im_out(22) => data_im_out(356),
            data_im_out(23) => data_im_out(372),
            data_im_out(24) => data_im_out(388),
            data_im_out(25) => data_im_out(404),
            data_im_out(26) => data_im_out(420),
            data_im_out(27) => data_im_out(436),
            data_im_out(28) => data_im_out(452),
            data_im_out(29) => data_im_out(468),
            data_im_out(30) => data_im_out(484),
            data_im_out(31) => data_im_out(500)
        );           

    URFFT_PT32_5 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(160),
            data_re_in(1) => mul_re_out(161),
            data_re_in(2) => mul_re_out(162),
            data_re_in(3) => mul_re_out(163),
            data_re_in(4) => mul_re_out(164),
            data_re_in(5) => mul_re_out(165),
            data_re_in(6) => mul_re_out(166),
            data_re_in(7) => mul_re_out(167),
            data_re_in(8) => mul_re_out(168),
            data_re_in(9) => mul_re_out(169),
            data_re_in(10) => mul_re_out(170),
            data_re_in(11) => mul_re_out(171),
            data_re_in(12) => mul_re_out(172),
            data_re_in(13) => mul_re_out(173),
            data_re_in(14) => mul_re_out(174),
            data_re_in(15) => mul_re_out(175),
            data_re_in(16) => mul_re_out(176),
            data_re_in(17) => mul_re_out(177),
            data_re_in(18) => mul_re_out(178),
            data_re_in(19) => mul_re_out(179),
            data_re_in(20) => mul_re_out(180),
            data_re_in(21) => mul_re_out(181),
            data_re_in(22) => mul_re_out(182),
            data_re_in(23) => mul_re_out(183),
            data_re_in(24) => mul_re_out(184),
            data_re_in(25) => mul_re_out(185),
            data_re_in(26) => mul_re_out(186),
            data_re_in(27) => mul_re_out(187),
            data_re_in(28) => mul_re_out(188),
            data_re_in(29) => mul_re_out(189),
            data_re_in(30) => mul_re_out(190),
            data_re_in(31) => mul_re_out(191),
            data_im_in(0) => mul_im_out(160),
            data_im_in(1) => mul_im_out(161),
            data_im_in(2) => mul_im_out(162),
            data_im_in(3) => mul_im_out(163),
            data_im_in(4) => mul_im_out(164),
            data_im_in(5) => mul_im_out(165),
            data_im_in(6) => mul_im_out(166),
            data_im_in(7) => mul_im_out(167),
            data_im_in(8) => mul_im_out(168),
            data_im_in(9) => mul_im_out(169),
            data_im_in(10) => mul_im_out(170),
            data_im_in(11) => mul_im_out(171),
            data_im_in(12) => mul_im_out(172),
            data_im_in(13) => mul_im_out(173),
            data_im_in(14) => mul_im_out(174),
            data_im_in(15) => mul_im_out(175),
            data_im_in(16) => mul_im_out(176),
            data_im_in(17) => mul_im_out(177),
            data_im_in(18) => mul_im_out(178),
            data_im_in(19) => mul_im_out(179),
            data_im_in(20) => mul_im_out(180),
            data_im_in(21) => mul_im_out(181),
            data_im_in(22) => mul_im_out(182),
            data_im_in(23) => mul_im_out(183),
            data_im_in(24) => mul_im_out(184),
            data_im_in(25) => mul_im_out(185),
            data_im_in(26) => mul_im_out(186),
            data_im_in(27) => mul_im_out(187),
            data_im_in(28) => mul_im_out(188),
            data_im_in(29) => mul_im_out(189),
            data_im_in(30) => mul_im_out(190),
            data_im_in(31) => mul_im_out(191),
            data_re_out(0) => data_re_out(5),
            data_re_out(1) => data_re_out(21),
            data_re_out(2) => data_re_out(37),
            data_re_out(3) => data_re_out(53),
            data_re_out(4) => data_re_out(69),
            data_re_out(5) => data_re_out(85),
            data_re_out(6) => data_re_out(101),
            data_re_out(7) => data_re_out(117),
            data_re_out(8) => data_re_out(133),
            data_re_out(9) => data_re_out(149),
            data_re_out(10) => data_re_out(165),
            data_re_out(11) => data_re_out(181),
            data_re_out(12) => data_re_out(197),
            data_re_out(13) => data_re_out(213),
            data_re_out(14) => data_re_out(229),
            data_re_out(15) => data_re_out(245),
            data_re_out(16) => data_re_out(261),
            data_re_out(17) => data_re_out(277),
            data_re_out(18) => data_re_out(293),
            data_re_out(19) => data_re_out(309),
            data_re_out(20) => data_re_out(325),
            data_re_out(21) => data_re_out(341),
            data_re_out(22) => data_re_out(357),
            data_re_out(23) => data_re_out(373),
            data_re_out(24) => data_re_out(389),
            data_re_out(25) => data_re_out(405),
            data_re_out(26) => data_re_out(421),
            data_re_out(27) => data_re_out(437),
            data_re_out(28) => data_re_out(453),
            data_re_out(29) => data_re_out(469),
            data_re_out(30) => data_re_out(485),
            data_re_out(31) => data_re_out(501),
            data_im_out(0) => data_im_out(5),
            data_im_out(1) => data_im_out(21),
            data_im_out(2) => data_im_out(37),
            data_im_out(3) => data_im_out(53),
            data_im_out(4) => data_im_out(69),
            data_im_out(5) => data_im_out(85),
            data_im_out(6) => data_im_out(101),
            data_im_out(7) => data_im_out(117),
            data_im_out(8) => data_im_out(133),
            data_im_out(9) => data_im_out(149),
            data_im_out(10) => data_im_out(165),
            data_im_out(11) => data_im_out(181),
            data_im_out(12) => data_im_out(197),
            data_im_out(13) => data_im_out(213),
            data_im_out(14) => data_im_out(229),
            data_im_out(15) => data_im_out(245),
            data_im_out(16) => data_im_out(261),
            data_im_out(17) => data_im_out(277),
            data_im_out(18) => data_im_out(293),
            data_im_out(19) => data_im_out(309),
            data_im_out(20) => data_im_out(325),
            data_im_out(21) => data_im_out(341),
            data_im_out(22) => data_im_out(357),
            data_im_out(23) => data_im_out(373),
            data_im_out(24) => data_im_out(389),
            data_im_out(25) => data_im_out(405),
            data_im_out(26) => data_im_out(421),
            data_im_out(27) => data_im_out(437),
            data_im_out(28) => data_im_out(453),
            data_im_out(29) => data_im_out(469),
            data_im_out(30) => data_im_out(485),
            data_im_out(31) => data_im_out(501)
        );           

    URFFT_PT32_6 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(192),
            data_re_in(1) => mul_re_out(193),
            data_re_in(2) => mul_re_out(194),
            data_re_in(3) => mul_re_out(195),
            data_re_in(4) => mul_re_out(196),
            data_re_in(5) => mul_re_out(197),
            data_re_in(6) => mul_re_out(198),
            data_re_in(7) => mul_re_out(199),
            data_re_in(8) => mul_re_out(200),
            data_re_in(9) => mul_re_out(201),
            data_re_in(10) => mul_re_out(202),
            data_re_in(11) => mul_re_out(203),
            data_re_in(12) => mul_re_out(204),
            data_re_in(13) => mul_re_out(205),
            data_re_in(14) => mul_re_out(206),
            data_re_in(15) => mul_re_out(207),
            data_re_in(16) => mul_re_out(208),
            data_re_in(17) => mul_re_out(209),
            data_re_in(18) => mul_re_out(210),
            data_re_in(19) => mul_re_out(211),
            data_re_in(20) => mul_re_out(212),
            data_re_in(21) => mul_re_out(213),
            data_re_in(22) => mul_re_out(214),
            data_re_in(23) => mul_re_out(215),
            data_re_in(24) => mul_re_out(216),
            data_re_in(25) => mul_re_out(217),
            data_re_in(26) => mul_re_out(218),
            data_re_in(27) => mul_re_out(219),
            data_re_in(28) => mul_re_out(220),
            data_re_in(29) => mul_re_out(221),
            data_re_in(30) => mul_re_out(222),
            data_re_in(31) => mul_re_out(223),
            data_im_in(0) => mul_im_out(192),
            data_im_in(1) => mul_im_out(193),
            data_im_in(2) => mul_im_out(194),
            data_im_in(3) => mul_im_out(195),
            data_im_in(4) => mul_im_out(196),
            data_im_in(5) => mul_im_out(197),
            data_im_in(6) => mul_im_out(198),
            data_im_in(7) => mul_im_out(199),
            data_im_in(8) => mul_im_out(200),
            data_im_in(9) => mul_im_out(201),
            data_im_in(10) => mul_im_out(202),
            data_im_in(11) => mul_im_out(203),
            data_im_in(12) => mul_im_out(204),
            data_im_in(13) => mul_im_out(205),
            data_im_in(14) => mul_im_out(206),
            data_im_in(15) => mul_im_out(207),
            data_im_in(16) => mul_im_out(208),
            data_im_in(17) => mul_im_out(209),
            data_im_in(18) => mul_im_out(210),
            data_im_in(19) => mul_im_out(211),
            data_im_in(20) => mul_im_out(212),
            data_im_in(21) => mul_im_out(213),
            data_im_in(22) => mul_im_out(214),
            data_im_in(23) => mul_im_out(215),
            data_im_in(24) => mul_im_out(216),
            data_im_in(25) => mul_im_out(217),
            data_im_in(26) => mul_im_out(218),
            data_im_in(27) => mul_im_out(219),
            data_im_in(28) => mul_im_out(220),
            data_im_in(29) => mul_im_out(221),
            data_im_in(30) => mul_im_out(222),
            data_im_in(31) => mul_im_out(223),
            data_re_out(0) => data_re_out(6),
            data_re_out(1) => data_re_out(22),
            data_re_out(2) => data_re_out(38),
            data_re_out(3) => data_re_out(54),
            data_re_out(4) => data_re_out(70),
            data_re_out(5) => data_re_out(86),
            data_re_out(6) => data_re_out(102),
            data_re_out(7) => data_re_out(118),
            data_re_out(8) => data_re_out(134),
            data_re_out(9) => data_re_out(150),
            data_re_out(10) => data_re_out(166),
            data_re_out(11) => data_re_out(182),
            data_re_out(12) => data_re_out(198),
            data_re_out(13) => data_re_out(214),
            data_re_out(14) => data_re_out(230),
            data_re_out(15) => data_re_out(246),
            data_re_out(16) => data_re_out(262),
            data_re_out(17) => data_re_out(278),
            data_re_out(18) => data_re_out(294),
            data_re_out(19) => data_re_out(310),
            data_re_out(20) => data_re_out(326),
            data_re_out(21) => data_re_out(342),
            data_re_out(22) => data_re_out(358),
            data_re_out(23) => data_re_out(374),
            data_re_out(24) => data_re_out(390),
            data_re_out(25) => data_re_out(406),
            data_re_out(26) => data_re_out(422),
            data_re_out(27) => data_re_out(438),
            data_re_out(28) => data_re_out(454),
            data_re_out(29) => data_re_out(470),
            data_re_out(30) => data_re_out(486),
            data_re_out(31) => data_re_out(502),
            data_im_out(0) => data_im_out(6),
            data_im_out(1) => data_im_out(22),
            data_im_out(2) => data_im_out(38),
            data_im_out(3) => data_im_out(54),
            data_im_out(4) => data_im_out(70),
            data_im_out(5) => data_im_out(86),
            data_im_out(6) => data_im_out(102),
            data_im_out(7) => data_im_out(118),
            data_im_out(8) => data_im_out(134),
            data_im_out(9) => data_im_out(150),
            data_im_out(10) => data_im_out(166),
            data_im_out(11) => data_im_out(182),
            data_im_out(12) => data_im_out(198),
            data_im_out(13) => data_im_out(214),
            data_im_out(14) => data_im_out(230),
            data_im_out(15) => data_im_out(246),
            data_im_out(16) => data_im_out(262),
            data_im_out(17) => data_im_out(278),
            data_im_out(18) => data_im_out(294),
            data_im_out(19) => data_im_out(310),
            data_im_out(20) => data_im_out(326),
            data_im_out(21) => data_im_out(342),
            data_im_out(22) => data_im_out(358),
            data_im_out(23) => data_im_out(374),
            data_im_out(24) => data_im_out(390),
            data_im_out(25) => data_im_out(406),
            data_im_out(26) => data_im_out(422),
            data_im_out(27) => data_im_out(438),
            data_im_out(28) => data_im_out(454),
            data_im_out(29) => data_im_out(470),
            data_im_out(30) => data_im_out(486),
            data_im_out(31) => data_im_out(502)
        );           

    URFFT_PT32_7 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(224),
            data_re_in(1) => mul_re_out(225),
            data_re_in(2) => mul_re_out(226),
            data_re_in(3) => mul_re_out(227),
            data_re_in(4) => mul_re_out(228),
            data_re_in(5) => mul_re_out(229),
            data_re_in(6) => mul_re_out(230),
            data_re_in(7) => mul_re_out(231),
            data_re_in(8) => mul_re_out(232),
            data_re_in(9) => mul_re_out(233),
            data_re_in(10) => mul_re_out(234),
            data_re_in(11) => mul_re_out(235),
            data_re_in(12) => mul_re_out(236),
            data_re_in(13) => mul_re_out(237),
            data_re_in(14) => mul_re_out(238),
            data_re_in(15) => mul_re_out(239),
            data_re_in(16) => mul_re_out(240),
            data_re_in(17) => mul_re_out(241),
            data_re_in(18) => mul_re_out(242),
            data_re_in(19) => mul_re_out(243),
            data_re_in(20) => mul_re_out(244),
            data_re_in(21) => mul_re_out(245),
            data_re_in(22) => mul_re_out(246),
            data_re_in(23) => mul_re_out(247),
            data_re_in(24) => mul_re_out(248),
            data_re_in(25) => mul_re_out(249),
            data_re_in(26) => mul_re_out(250),
            data_re_in(27) => mul_re_out(251),
            data_re_in(28) => mul_re_out(252),
            data_re_in(29) => mul_re_out(253),
            data_re_in(30) => mul_re_out(254),
            data_re_in(31) => mul_re_out(255),
            data_im_in(0) => mul_im_out(224),
            data_im_in(1) => mul_im_out(225),
            data_im_in(2) => mul_im_out(226),
            data_im_in(3) => mul_im_out(227),
            data_im_in(4) => mul_im_out(228),
            data_im_in(5) => mul_im_out(229),
            data_im_in(6) => mul_im_out(230),
            data_im_in(7) => mul_im_out(231),
            data_im_in(8) => mul_im_out(232),
            data_im_in(9) => mul_im_out(233),
            data_im_in(10) => mul_im_out(234),
            data_im_in(11) => mul_im_out(235),
            data_im_in(12) => mul_im_out(236),
            data_im_in(13) => mul_im_out(237),
            data_im_in(14) => mul_im_out(238),
            data_im_in(15) => mul_im_out(239),
            data_im_in(16) => mul_im_out(240),
            data_im_in(17) => mul_im_out(241),
            data_im_in(18) => mul_im_out(242),
            data_im_in(19) => mul_im_out(243),
            data_im_in(20) => mul_im_out(244),
            data_im_in(21) => mul_im_out(245),
            data_im_in(22) => mul_im_out(246),
            data_im_in(23) => mul_im_out(247),
            data_im_in(24) => mul_im_out(248),
            data_im_in(25) => mul_im_out(249),
            data_im_in(26) => mul_im_out(250),
            data_im_in(27) => mul_im_out(251),
            data_im_in(28) => mul_im_out(252),
            data_im_in(29) => mul_im_out(253),
            data_im_in(30) => mul_im_out(254),
            data_im_in(31) => mul_im_out(255),
            data_re_out(0) => data_re_out(7),
            data_re_out(1) => data_re_out(23),
            data_re_out(2) => data_re_out(39),
            data_re_out(3) => data_re_out(55),
            data_re_out(4) => data_re_out(71),
            data_re_out(5) => data_re_out(87),
            data_re_out(6) => data_re_out(103),
            data_re_out(7) => data_re_out(119),
            data_re_out(8) => data_re_out(135),
            data_re_out(9) => data_re_out(151),
            data_re_out(10) => data_re_out(167),
            data_re_out(11) => data_re_out(183),
            data_re_out(12) => data_re_out(199),
            data_re_out(13) => data_re_out(215),
            data_re_out(14) => data_re_out(231),
            data_re_out(15) => data_re_out(247),
            data_re_out(16) => data_re_out(263),
            data_re_out(17) => data_re_out(279),
            data_re_out(18) => data_re_out(295),
            data_re_out(19) => data_re_out(311),
            data_re_out(20) => data_re_out(327),
            data_re_out(21) => data_re_out(343),
            data_re_out(22) => data_re_out(359),
            data_re_out(23) => data_re_out(375),
            data_re_out(24) => data_re_out(391),
            data_re_out(25) => data_re_out(407),
            data_re_out(26) => data_re_out(423),
            data_re_out(27) => data_re_out(439),
            data_re_out(28) => data_re_out(455),
            data_re_out(29) => data_re_out(471),
            data_re_out(30) => data_re_out(487),
            data_re_out(31) => data_re_out(503),
            data_im_out(0) => data_im_out(7),
            data_im_out(1) => data_im_out(23),
            data_im_out(2) => data_im_out(39),
            data_im_out(3) => data_im_out(55),
            data_im_out(4) => data_im_out(71),
            data_im_out(5) => data_im_out(87),
            data_im_out(6) => data_im_out(103),
            data_im_out(7) => data_im_out(119),
            data_im_out(8) => data_im_out(135),
            data_im_out(9) => data_im_out(151),
            data_im_out(10) => data_im_out(167),
            data_im_out(11) => data_im_out(183),
            data_im_out(12) => data_im_out(199),
            data_im_out(13) => data_im_out(215),
            data_im_out(14) => data_im_out(231),
            data_im_out(15) => data_im_out(247),
            data_im_out(16) => data_im_out(263),
            data_im_out(17) => data_im_out(279),
            data_im_out(18) => data_im_out(295),
            data_im_out(19) => data_im_out(311),
            data_im_out(20) => data_im_out(327),
            data_im_out(21) => data_im_out(343),
            data_im_out(22) => data_im_out(359),
            data_im_out(23) => data_im_out(375),
            data_im_out(24) => data_im_out(391),
            data_im_out(25) => data_im_out(407),
            data_im_out(26) => data_im_out(423),
            data_im_out(27) => data_im_out(439),
            data_im_out(28) => data_im_out(455),
            data_im_out(29) => data_im_out(471),
            data_im_out(30) => data_im_out(487),
            data_im_out(31) => data_im_out(503)
        );           

    URFFT_PT32_8 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(256),
            data_re_in(1) => mul_re_out(257),
            data_re_in(2) => mul_re_out(258),
            data_re_in(3) => mul_re_out(259),
            data_re_in(4) => mul_re_out(260),
            data_re_in(5) => mul_re_out(261),
            data_re_in(6) => mul_re_out(262),
            data_re_in(7) => mul_re_out(263),
            data_re_in(8) => mul_re_out(264),
            data_re_in(9) => mul_re_out(265),
            data_re_in(10) => mul_re_out(266),
            data_re_in(11) => mul_re_out(267),
            data_re_in(12) => mul_re_out(268),
            data_re_in(13) => mul_re_out(269),
            data_re_in(14) => mul_re_out(270),
            data_re_in(15) => mul_re_out(271),
            data_re_in(16) => mul_re_out(272),
            data_re_in(17) => mul_re_out(273),
            data_re_in(18) => mul_re_out(274),
            data_re_in(19) => mul_re_out(275),
            data_re_in(20) => mul_re_out(276),
            data_re_in(21) => mul_re_out(277),
            data_re_in(22) => mul_re_out(278),
            data_re_in(23) => mul_re_out(279),
            data_re_in(24) => mul_re_out(280),
            data_re_in(25) => mul_re_out(281),
            data_re_in(26) => mul_re_out(282),
            data_re_in(27) => mul_re_out(283),
            data_re_in(28) => mul_re_out(284),
            data_re_in(29) => mul_re_out(285),
            data_re_in(30) => mul_re_out(286),
            data_re_in(31) => mul_re_out(287),
            data_im_in(0) => mul_im_out(256),
            data_im_in(1) => mul_im_out(257),
            data_im_in(2) => mul_im_out(258),
            data_im_in(3) => mul_im_out(259),
            data_im_in(4) => mul_im_out(260),
            data_im_in(5) => mul_im_out(261),
            data_im_in(6) => mul_im_out(262),
            data_im_in(7) => mul_im_out(263),
            data_im_in(8) => mul_im_out(264),
            data_im_in(9) => mul_im_out(265),
            data_im_in(10) => mul_im_out(266),
            data_im_in(11) => mul_im_out(267),
            data_im_in(12) => mul_im_out(268),
            data_im_in(13) => mul_im_out(269),
            data_im_in(14) => mul_im_out(270),
            data_im_in(15) => mul_im_out(271),
            data_im_in(16) => mul_im_out(272),
            data_im_in(17) => mul_im_out(273),
            data_im_in(18) => mul_im_out(274),
            data_im_in(19) => mul_im_out(275),
            data_im_in(20) => mul_im_out(276),
            data_im_in(21) => mul_im_out(277),
            data_im_in(22) => mul_im_out(278),
            data_im_in(23) => mul_im_out(279),
            data_im_in(24) => mul_im_out(280),
            data_im_in(25) => mul_im_out(281),
            data_im_in(26) => mul_im_out(282),
            data_im_in(27) => mul_im_out(283),
            data_im_in(28) => mul_im_out(284),
            data_im_in(29) => mul_im_out(285),
            data_im_in(30) => mul_im_out(286),
            data_im_in(31) => mul_im_out(287),
            data_re_out(0) => data_re_out(8),
            data_re_out(1) => data_re_out(24),
            data_re_out(2) => data_re_out(40),
            data_re_out(3) => data_re_out(56),
            data_re_out(4) => data_re_out(72),
            data_re_out(5) => data_re_out(88),
            data_re_out(6) => data_re_out(104),
            data_re_out(7) => data_re_out(120),
            data_re_out(8) => data_re_out(136),
            data_re_out(9) => data_re_out(152),
            data_re_out(10) => data_re_out(168),
            data_re_out(11) => data_re_out(184),
            data_re_out(12) => data_re_out(200),
            data_re_out(13) => data_re_out(216),
            data_re_out(14) => data_re_out(232),
            data_re_out(15) => data_re_out(248),
            data_re_out(16) => data_re_out(264),
            data_re_out(17) => data_re_out(280),
            data_re_out(18) => data_re_out(296),
            data_re_out(19) => data_re_out(312),
            data_re_out(20) => data_re_out(328),
            data_re_out(21) => data_re_out(344),
            data_re_out(22) => data_re_out(360),
            data_re_out(23) => data_re_out(376),
            data_re_out(24) => data_re_out(392),
            data_re_out(25) => data_re_out(408),
            data_re_out(26) => data_re_out(424),
            data_re_out(27) => data_re_out(440),
            data_re_out(28) => data_re_out(456),
            data_re_out(29) => data_re_out(472),
            data_re_out(30) => data_re_out(488),
            data_re_out(31) => data_re_out(504),
            data_im_out(0) => data_im_out(8),
            data_im_out(1) => data_im_out(24),
            data_im_out(2) => data_im_out(40),
            data_im_out(3) => data_im_out(56),
            data_im_out(4) => data_im_out(72),
            data_im_out(5) => data_im_out(88),
            data_im_out(6) => data_im_out(104),
            data_im_out(7) => data_im_out(120),
            data_im_out(8) => data_im_out(136),
            data_im_out(9) => data_im_out(152),
            data_im_out(10) => data_im_out(168),
            data_im_out(11) => data_im_out(184),
            data_im_out(12) => data_im_out(200),
            data_im_out(13) => data_im_out(216),
            data_im_out(14) => data_im_out(232),
            data_im_out(15) => data_im_out(248),
            data_im_out(16) => data_im_out(264),
            data_im_out(17) => data_im_out(280),
            data_im_out(18) => data_im_out(296),
            data_im_out(19) => data_im_out(312),
            data_im_out(20) => data_im_out(328),
            data_im_out(21) => data_im_out(344),
            data_im_out(22) => data_im_out(360),
            data_im_out(23) => data_im_out(376),
            data_im_out(24) => data_im_out(392),
            data_im_out(25) => data_im_out(408),
            data_im_out(26) => data_im_out(424),
            data_im_out(27) => data_im_out(440),
            data_im_out(28) => data_im_out(456),
            data_im_out(29) => data_im_out(472),
            data_im_out(30) => data_im_out(488),
            data_im_out(31) => data_im_out(504)
        );           

    URFFT_PT32_9 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(288),
            data_re_in(1) => mul_re_out(289),
            data_re_in(2) => mul_re_out(290),
            data_re_in(3) => mul_re_out(291),
            data_re_in(4) => mul_re_out(292),
            data_re_in(5) => mul_re_out(293),
            data_re_in(6) => mul_re_out(294),
            data_re_in(7) => mul_re_out(295),
            data_re_in(8) => mul_re_out(296),
            data_re_in(9) => mul_re_out(297),
            data_re_in(10) => mul_re_out(298),
            data_re_in(11) => mul_re_out(299),
            data_re_in(12) => mul_re_out(300),
            data_re_in(13) => mul_re_out(301),
            data_re_in(14) => mul_re_out(302),
            data_re_in(15) => mul_re_out(303),
            data_re_in(16) => mul_re_out(304),
            data_re_in(17) => mul_re_out(305),
            data_re_in(18) => mul_re_out(306),
            data_re_in(19) => mul_re_out(307),
            data_re_in(20) => mul_re_out(308),
            data_re_in(21) => mul_re_out(309),
            data_re_in(22) => mul_re_out(310),
            data_re_in(23) => mul_re_out(311),
            data_re_in(24) => mul_re_out(312),
            data_re_in(25) => mul_re_out(313),
            data_re_in(26) => mul_re_out(314),
            data_re_in(27) => mul_re_out(315),
            data_re_in(28) => mul_re_out(316),
            data_re_in(29) => mul_re_out(317),
            data_re_in(30) => mul_re_out(318),
            data_re_in(31) => mul_re_out(319),
            data_im_in(0) => mul_im_out(288),
            data_im_in(1) => mul_im_out(289),
            data_im_in(2) => mul_im_out(290),
            data_im_in(3) => mul_im_out(291),
            data_im_in(4) => mul_im_out(292),
            data_im_in(5) => mul_im_out(293),
            data_im_in(6) => mul_im_out(294),
            data_im_in(7) => mul_im_out(295),
            data_im_in(8) => mul_im_out(296),
            data_im_in(9) => mul_im_out(297),
            data_im_in(10) => mul_im_out(298),
            data_im_in(11) => mul_im_out(299),
            data_im_in(12) => mul_im_out(300),
            data_im_in(13) => mul_im_out(301),
            data_im_in(14) => mul_im_out(302),
            data_im_in(15) => mul_im_out(303),
            data_im_in(16) => mul_im_out(304),
            data_im_in(17) => mul_im_out(305),
            data_im_in(18) => mul_im_out(306),
            data_im_in(19) => mul_im_out(307),
            data_im_in(20) => mul_im_out(308),
            data_im_in(21) => mul_im_out(309),
            data_im_in(22) => mul_im_out(310),
            data_im_in(23) => mul_im_out(311),
            data_im_in(24) => mul_im_out(312),
            data_im_in(25) => mul_im_out(313),
            data_im_in(26) => mul_im_out(314),
            data_im_in(27) => mul_im_out(315),
            data_im_in(28) => mul_im_out(316),
            data_im_in(29) => mul_im_out(317),
            data_im_in(30) => mul_im_out(318),
            data_im_in(31) => mul_im_out(319),
            data_re_out(0) => data_re_out(9),
            data_re_out(1) => data_re_out(25),
            data_re_out(2) => data_re_out(41),
            data_re_out(3) => data_re_out(57),
            data_re_out(4) => data_re_out(73),
            data_re_out(5) => data_re_out(89),
            data_re_out(6) => data_re_out(105),
            data_re_out(7) => data_re_out(121),
            data_re_out(8) => data_re_out(137),
            data_re_out(9) => data_re_out(153),
            data_re_out(10) => data_re_out(169),
            data_re_out(11) => data_re_out(185),
            data_re_out(12) => data_re_out(201),
            data_re_out(13) => data_re_out(217),
            data_re_out(14) => data_re_out(233),
            data_re_out(15) => data_re_out(249),
            data_re_out(16) => data_re_out(265),
            data_re_out(17) => data_re_out(281),
            data_re_out(18) => data_re_out(297),
            data_re_out(19) => data_re_out(313),
            data_re_out(20) => data_re_out(329),
            data_re_out(21) => data_re_out(345),
            data_re_out(22) => data_re_out(361),
            data_re_out(23) => data_re_out(377),
            data_re_out(24) => data_re_out(393),
            data_re_out(25) => data_re_out(409),
            data_re_out(26) => data_re_out(425),
            data_re_out(27) => data_re_out(441),
            data_re_out(28) => data_re_out(457),
            data_re_out(29) => data_re_out(473),
            data_re_out(30) => data_re_out(489),
            data_re_out(31) => data_re_out(505),
            data_im_out(0) => data_im_out(9),
            data_im_out(1) => data_im_out(25),
            data_im_out(2) => data_im_out(41),
            data_im_out(3) => data_im_out(57),
            data_im_out(4) => data_im_out(73),
            data_im_out(5) => data_im_out(89),
            data_im_out(6) => data_im_out(105),
            data_im_out(7) => data_im_out(121),
            data_im_out(8) => data_im_out(137),
            data_im_out(9) => data_im_out(153),
            data_im_out(10) => data_im_out(169),
            data_im_out(11) => data_im_out(185),
            data_im_out(12) => data_im_out(201),
            data_im_out(13) => data_im_out(217),
            data_im_out(14) => data_im_out(233),
            data_im_out(15) => data_im_out(249),
            data_im_out(16) => data_im_out(265),
            data_im_out(17) => data_im_out(281),
            data_im_out(18) => data_im_out(297),
            data_im_out(19) => data_im_out(313),
            data_im_out(20) => data_im_out(329),
            data_im_out(21) => data_im_out(345),
            data_im_out(22) => data_im_out(361),
            data_im_out(23) => data_im_out(377),
            data_im_out(24) => data_im_out(393),
            data_im_out(25) => data_im_out(409),
            data_im_out(26) => data_im_out(425),
            data_im_out(27) => data_im_out(441),
            data_im_out(28) => data_im_out(457),
            data_im_out(29) => data_im_out(473),
            data_im_out(30) => data_im_out(489),
            data_im_out(31) => data_im_out(505)
        );           

    URFFT_PT32_10 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(320),
            data_re_in(1) => mul_re_out(321),
            data_re_in(2) => mul_re_out(322),
            data_re_in(3) => mul_re_out(323),
            data_re_in(4) => mul_re_out(324),
            data_re_in(5) => mul_re_out(325),
            data_re_in(6) => mul_re_out(326),
            data_re_in(7) => mul_re_out(327),
            data_re_in(8) => mul_re_out(328),
            data_re_in(9) => mul_re_out(329),
            data_re_in(10) => mul_re_out(330),
            data_re_in(11) => mul_re_out(331),
            data_re_in(12) => mul_re_out(332),
            data_re_in(13) => mul_re_out(333),
            data_re_in(14) => mul_re_out(334),
            data_re_in(15) => mul_re_out(335),
            data_re_in(16) => mul_re_out(336),
            data_re_in(17) => mul_re_out(337),
            data_re_in(18) => mul_re_out(338),
            data_re_in(19) => mul_re_out(339),
            data_re_in(20) => mul_re_out(340),
            data_re_in(21) => mul_re_out(341),
            data_re_in(22) => mul_re_out(342),
            data_re_in(23) => mul_re_out(343),
            data_re_in(24) => mul_re_out(344),
            data_re_in(25) => mul_re_out(345),
            data_re_in(26) => mul_re_out(346),
            data_re_in(27) => mul_re_out(347),
            data_re_in(28) => mul_re_out(348),
            data_re_in(29) => mul_re_out(349),
            data_re_in(30) => mul_re_out(350),
            data_re_in(31) => mul_re_out(351),
            data_im_in(0) => mul_im_out(320),
            data_im_in(1) => mul_im_out(321),
            data_im_in(2) => mul_im_out(322),
            data_im_in(3) => mul_im_out(323),
            data_im_in(4) => mul_im_out(324),
            data_im_in(5) => mul_im_out(325),
            data_im_in(6) => mul_im_out(326),
            data_im_in(7) => mul_im_out(327),
            data_im_in(8) => mul_im_out(328),
            data_im_in(9) => mul_im_out(329),
            data_im_in(10) => mul_im_out(330),
            data_im_in(11) => mul_im_out(331),
            data_im_in(12) => mul_im_out(332),
            data_im_in(13) => mul_im_out(333),
            data_im_in(14) => mul_im_out(334),
            data_im_in(15) => mul_im_out(335),
            data_im_in(16) => mul_im_out(336),
            data_im_in(17) => mul_im_out(337),
            data_im_in(18) => mul_im_out(338),
            data_im_in(19) => mul_im_out(339),
            data_im_in(20) => mul_im_out(340),
            data_im_in(21) => mul_im_out(341),
            data_im_in(22) => mul_im_out(342),
            data_im_in(23) => mul_im_out(343),
            data_im_in(24) => mul_im_out(344),
            data_im_in(25) => mul_im_out(345),
            data_im_in(26) => mul_im_out(346),
            data_im_in(27) => mul_im_out(347),
            data_im_in(28) => mul_im_out(348),
            data_im_in(29) => mul_im_out(349),
            data_im_in(30) => mul_im_out(350),
            data_im_in(31) => mul_im_out(351),
            data_re_out(0) => data_re_out(10),
            data_re_out(1) => data_re_out(26),
            data_re_out(2) => data_re_out(42),
            data_re_out(3) => data_re_out(58),
            data_re_out(4) => data_re_out(74),
            data_re_out(5) => data_re_out(90),
            data_re_out(6) => data_re_out(106),
            data_re_out(7) => data_re_out(122),
            data_re_out(8) => data_re_out(138),
            data_re_out(9) => data_re_out(154),
            data_re_out(10) => data_re_out(170),
            data_re_out(11) => data_re_out(186),
            data_re_out(12) => data_re_out(202),
            data_re_out(13) => data_re_out(218),
            data_re_out(14) => data_re_out(234),
            data_re_out(15) => data_re_out(250),
            data_re_out(16) => data_re_out(266),
            data_re_out(17) => data_re_out(282),
            data_re_out(18) => data_re_out(298),
            data_re_out(19) => data_re_out(314),
            data_re_out(20) => data_re_out(330),
            data_re_out(21) => data_re_out(346),
            data_re_out(22) => data_re_out(362),
            data_re_out(23) => data_re_out(378),
            data_re_out(24) => data_re_out(394),
            data_re_out(25) => data_re_out(410),
            data_re_out(26) => data_re_out(426),
            data_re_out(27) => data_re_out(442),
            data_re_out(28) => data_re_out(458),
            data_re_out(29) => data_re_out(474),
            data_re_out(30) => data_re_out(490),
            data_re_out(31) => data_re_out(506),
            data_im_out(0) => data_im_out(10),
            data_im_out(1) => data_im_out(26),
            data_im_out(2) => data_im_out(42),
            data_im_out(3) => data_im_out(58),
            data_im_out(4) => data_im_out(74),
            data_im_out(5) => data_im_out(90),
            data_im_out(6) => data_im_out(106),
            data_im_out(7) => data_im_out(122),
            data_im_out(8) => data_im_out(138),
            data_im_out(9) => data_im_out(154),
            data_im_out(10) => data_im_out(170),
            data_im_out(11) => data_im_out(186),
            data_im_out(12) => data_im_out(202),
            data_im_out(13) => data_im_out(218),
            data_im_out(14) => data_im_out(234),
            data_im_out(15) => data_im_out(250),
            data_im_out(16) => data_im_out(266),
            data_im_out(17) => data_im_out(282),
            data_im_out(18) => data_im_out(298),
            data_im_out(19) => data_im_out(314),
            data_im_out(20) => data_im_out(330),
            data_im_out(21) => data_im_out(346),
            data_im_out(22) => data_im_out(362),
            data_im_out(23) => data_im_out(378),
            data_im_out(24) => data_im_out(394),
            data_im_out(25) => data_im_out(410),
            data_im_out(26) => data_im_out(426),
            data_im_out(27) => data_im_out(442),
            data_im_out(28) => data_im_out(458),
            data_im_out(29) => data_im_out(474),
            data_im_out(30) => data_im_out(490),
            data_im_out(31) => data_im_out(506)
        );           

    URFFT_PT32_11 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(352),
            data_re_in(1) => mul_re_out(353),
            data_re_in(2) => mul_re_out(354),
            data_re_in(3) => mul_re_out(355),
            data_re_in(4) => mul_re_out(356),
            data_re_in(5) => mul_re_out(357),
            data_re_in(6) => mul_re_out(358),
            data_re_in(7) => mul_re_out(359),
            data_re_in(8) => mul_re_out(360),
            data_re_in(9) => mul_re_out(361),
            data_re_in(10) => mul_re_out(362),
            data_re_in(11) => mul_re_out(363),
            data_re_in(12) => mul_re_out(364),
            data_re_in(13) => mul_re_out(365),
            data_re_in(14) => mul_re_out(366),
            data_re_in(15) => mul_re_out(367),
            data_re_in(16) => mul_re_out(368),
            data_re_in(17) => mul_re_out(369),
            data_re_in(18) => mul_re_out(370),
            data_re_in(19) => mul_re_out(371),
            data_re_in(20) => mul_re_out(372),
            data_re_in(21) => mul_re_out(373),
            data_re_in(22) => mul_re_out(374),
            data_re_in(23) => mul_re_out(375),
            data_re_in(24) => mul_re_out(376),
            data_re_in(25) => mul_re_out(377),
            data_re_in(26) => mul_re_out(378),
            data_re_in(27) => mul_re_out(379),
            data_re_in(28) => mul_re_out(380),
            data_re_in(29) => mul_re_out(381),
            data_re_in(30) => mul_re_out(382),
            data_re_in(31) => mul_re_out(383),
            data_im_in(0) => mul_im_out(352),
            data_im_in(1) => mul_im_out(353),
            data_im_in(2) => mul_im_out(354),
            data_im_in(3) => mul_im_out(355),
            data_im_in(4) => mul_im_out(356),
            data_im_in(5) => mul_im_out(357),
            data_im_in(6) => mul_im_out(358),
            data_im_in(7) => mul_im_out(359),
            data_im_in(8) => mul_im_out(360),
            data_im_in(9) => mul_im_out(361),
            data_im_in(10) => mul_im_out(362),
            data_im_in(11) => mul_im_out(363),
            data_im_in(12) => mul_im_out(364),
            data_im_in(13) => mul_im_out(365),
            data_im_in(14) => mul_im_out(366),
            data_im_in(15) => mul_im_out(367),
            data_im_in(16) => mul_im_out(368),
            data_im_in(17) => mul_im_out(369),
            data_im_in(18) => mul_im_out(370),
            data_im_in(19) => mul_im_out(371),
            data_im_in(20) => mul_im_out(372),
            data_im_in(21) => mul_im_out(373),
            data_im_in(22) => mul_im_out(374),
            data_im_in(23) => mul_im_out(375),
            data_im_in(24) => mul_im_out(376),
            data_im_in(25) => mul_im_out(377),
            data_im_in(26) => mul_im_out(378),
            data_im_in(27) => mul_im_out(379),
            data_im_in(28) => mul_im_out(380),
            data_im_in(29) => mul_im_out(381),
            data_im_in(30) => mul_im_out(382),
            data_im_in(31) => mul_im_out(383),
            data_re_out(0) => data_re_out(11),
            data_re_out(1) => data_re_out(27),
            data_re_out(2) => data_re_out(43),
            data_re_out(3) => data_re_out(59),
            data_re_out(4) => data_re_out(75),
            data_re_out(5) => data_re_out(91),
            data_re_out(6) => data_re_out(107),
            data_re_out(7) => data_re_out(123),
            data_re_out(8) => data_re_out(139),
            data_re_out(9) => data_re_out(155),
            data_re_out(10) => data_re_out(171),
            data_re_out(11) => data_re_out(187),
            data_re_out(12) => data_re_out(203),
            data_re_out(13) => data_re_out(219),
            data_re_out(14) => data_re_out(235),
            data_re_out(15) => data_re_out(251),
            data_re_out(16) => data_re_out(267),
            data_re_out(17) => data_re_out(283),
            data_re_out(18) => data_re_out(299),
            data_re_out(19) => data_re_out(315),
            data_re_out(20) => data_re_out(331),
            data_re_out(21) => data_re_out(347),
            data_re_out(22) => data_re_out(363),
            data_re_out(23) => data_re_out(379),
            data_re_out(24) => data_re_out(395),
            data_re_out(25) => data_re_out(411),
            data_re_out(26) => data_re_out(427),
            data_re_out(27) => data_re_out(443),
            data_re_out(28) => data_re_out(459),
            data_re_out(29) => data_re_out(475),
            data_re_out(30) => data_re_out(491),
            data_re_out(31) => data_re_out(507),
            data_im_out(0) => data_im_out(11),
            data_im_out(1) => data_im_out(27),
            data_im_out(2) => data_im_out(43),
            data_im_out(3) => data_im_out(59),
            data_im_out(4) => data_im_out(75),
            data_im_out(5) => data_im_out(91),
            data_im_out(6) => data_im_out(107),
            data_im_out(7) => data_im_out(123),
            data_im_out(8) => data_im_out(139),
            data_im_out(9) => data_im_out(155),
            data_im_out(10) => data_im_out(171),
            data_im_out(11) => data_im_out(187),
            data_im_out(12) => data_im_out(203),
            data_im_out(13) => data_im_out(219),
            data_im_out(14) => data_im_out(235),
            data_im_out(15) => data_im_out(251),
            data_im_out(16) => data_im_out(267),
            data_im_out(17) => data_im_out(283),
            data_im_out(18) => data_im_out(299),
            data_im_out(19) => data_im_out(315),
            data_im_out(20) => data_im_out(331),
            data_im_out(21) => data_im_out(347),
            data_im_out(22) => data_im_out(363),
            data_im_out(23) => data_im_out(379),
            data_im_out(24) => data_im_out(395),
            data_im_out(25) => data_im_out(411),
            data_im_out(26) => data_im_out(427),
            data_im_out(27) => data_im_out(443),
            data_im_out(28) => data_im_out(459),
            data_im_out(29) => data_im_out(475),
            data_im_out(30) => data_im_out(491),
            data_im_out(31) => data_im_out(507)
        );           

    URFFT_PT32_12 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(384),
            data_re_in(1) => mul_re_out(385),
            data_re_in(2) => mul_re_out(386),
            data_re_in(3) => mul_re_out(387),
            data_re_in(4) => mul_re_out(388),
            data_re_in(5) => mul_re_out(389),
            data_re_in(6) => mul_re_out(390),
            data_re_in(7) => mul_re_out(391),
            data_re_in(8) => mul_re_out(392),
            data_re_in(9) => mul_re_out(393),
            data_re_in(10) => mul_re_out(394),
            data_re_in(11) => mul_re_out(395),
            data_re_in(12) => mul_re_out(396),
            data_re_in(13) => mul_re_out(397),
            data_re_in(14) => mul_re_out(398),
            data_re_in(15) => mul_re_out(399),
            data_re_in(16) => mul_re_out(400),
            data_re_in(17) => mul_re_out(401),
            data_re_in(18) => mul_re_out(402),
            data_re_in(19) => mul_re_out(403),
            data_re_in(20) => mul_re_out(404),
            data_re_in(21) => mul_re_out(405),
            data_re_in(22) => mul_re_out(406),
            data_re_in(23) => mul_re_out(407),
            data_re_in(24) => mul_re_out(408),
            data_re_in(25) => mul_re_out(409),
            data_re_in(26) => mul_re_out(410),
            data_re_in(27) => mul_re_out(411),
            data_re_in(28) => mul_re_out(412),
            data_re_in(29) => mul_re_out(413),
            data_re_in(30) => mul_re_out(414),
            data_re_in(31) => mul_re_out(415),
            data_im_in(0) => mul_im_out(384),
            data_im_in(1) => mul_im_out(385),
            data_im_in(2) => mul_im_out(386),
            data_im_in(3) => mul_im_out(387),
            data_im_in(4) => mul_im_out(388),
            data_im_in(5) => mul_im_out(389),
            data_im_in(6) => mul_im_out(390),
            data_im_in(7) => mul_im_out(391),
            data_im_in(8) => mul_im_out(392),
            data_im_in(9) => mul_im_out(393),
            data_im_in(10) => mul_im_out(394),
            data_im_in(11) => mul_im_out(395),
            data_im_in(12) => mul_im_out(396),
            data_im_in(13) => mul_im_out(397),
            data_im_in(14) => mul_im_out(398),
            data_im_in(15) => mul_im_out(399),
            data_im_in(16) => mul_im_out(400),
            data_im_in(17) => mul_im_out(401),
            data_im_in(18) => mul_im_out(402),
            data_im_in(19) => mul_im_out(403),
            data_im_in(20) => mul_im_out(404),
            data_im_in(21) => mul_im_out(405),
            data_im_in(22) => mul_im_out(406),
            data_im_in(23) => mul_im_out(407),
            data_im_in(24) => mul_im_out(408),
            data_im_in(25) => mul_im_out(409),
            data_im_in(26) => mul_im_out(410),
            data_im_in(27) => mul_im_out(411),
            data_im_in(28) => mul_im_out(412),
            data_im_in(29) => mul_im_out(413),
            data_im_in(30) => mul_im_out(414),
            data_im_in(31) => mul_im_out(415),
            data_re_out(0) => data_re_out(12),
            data_re_out(1) => data_re_out(28),
            data_re_out(2) => data_re_out(44),
            data_re_out(3) => data_re_out(60),
            data_re_out(4) => data_re_out(76),
            data_re_out(5) => data_re_out(92),
            data_re_out(6) => data_re_out(108),
            data_re_out(7) => data_re_out(124),
            data_re_out(8) => data_re_out(140),
            data_re_out(9) => data_re_out(156),
            data_re_out(10) => data_re_out(172),
            data_re_out(11) => data_re_out(188),
            data_re_out(12) => data_re_out(204),
            data_re_out(13) => data_re_out(220),
            data_re_out(14) => data_re_out(236),
            data_re_out(15) => data_re_out(252),
            data_re_out(16) => data_re_out(268),
            data_re_out(17) => data_re_out(284),
            data_re_out(18) => data_re_out(300),
            data_re_out(19) => data_re_out(316),
            data_re_out(20) => data_re_out(332),
            data_re_out(21) => data_re_out(348),
            data_re_out(22) => data_re_out(364),
            data_re_out(23) => data_re_out(380),
            data_re_out(24) => data_re_out(396),
            data_re_out(25) => data_re_out(412),
            data_re_out(26) => data_re_out(428),
            data_re_out(27) => data_re_out(444),
            data_re_out(28) => data_re_out(460),
            data_re_out(29) => data_re_out(476),
            data_re_out(30) => data_re_out(492),
            data_re_out(31) => data_re_out(508),
            data_im_out(0) => data_im_out(12),
            data_im_out(1) => data_im_out(28),
            data_im_out(2) => data_im_out(44),
            data_im_out(3) => data_im_out(60),
            data_im_out(4) => data_im_out(76),
            data_im_out(5) => data_im_out(92),
            data_im_out(6) => data_im_out(108),
            data_im_out(7) => data_im_out(124),
            data_im_out(8) => data_im_out(140),
            data_im_out(9) => data_im_out(156),
            data_im_out(10) => data_im_out(172),
            data_im_out(11) => data_im_out(188),
            data_im_out(12) => data_im_out(204),
            data_im_out(13) => data_im_out(220),
            data_im_out(14) => data_im_out(236),
            data_im_out(15) => data_im_out(252),
            data_im_out(16) => data_im_out(268),
            data_im_out(17) => data_im_out(284),
            data_im_out(18) => data_im_out(300),
            data_im_out(19) => data_im_out(316),
            data_im_out(20) => data_im_out(332),
            data_im_out(21) => data_im_out(348),
            data_im_out(22) => data_im_out(364),
            data_im_out(23) => data_im_out(380),
            data_im_out(24) => data_im_out(396),
            data_im_out(25) => data_im_out(412),
            data_im_out(26) => data_im_out(428),
            data_im_out(27) => data_im_out(444),
            data_im_out(28) => data_im_out(460),
            data_im_out(29) => data_im_out(476),
            data_im_out(30) => data_im_out(492),
            data_im_out(31) => data_im_out(508)
        );           

    URFFT_PT32_13 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(416),
            data_re_in(1) => mul_re_out(417),
            data_re_in(2) => mul_re_out(418),
            data_re_in(3) => mul_re_out(419),
            data_re_in(4) => mul_re_out(420),
            data_re_in(5) => mul_re_out(421),
            data_re_in(6) => mul_re_out(422),
            data_re_in(7) => mul_re_out(423),
            data_re_in(8) => mul_re_out(424),
            data_re_in(9) => mul_re_out(425),
            data_re_in(10) => mul_re_out(426),
            data_re_in(11) => mul_re_out(427),
            data_re_in(12) => mul_re_out(428),
            data_re_in(13) => mul_re_out(429),
            data_re_in(14) => mul_re_out(430),
            data_re_in(15) => mul_re_out(431),
            data_re_in(16) => mul_re_out(432),
            data_re_in(17) => mul_re_out(433),
            data_re_in(18) => mul_re_out(434),
            data_re_in(19) => mul_re_out(435),
            data_re_in(20) => mul_re_out(436),
            data_re_in(21) => mul_re_out(437),
            data_re_in(22) => mul_re_out(438),
            data_re_in(23) => mul_re_out(439),
            data_re_in(24) => mul_re_out(440),
            data_re_in(25) => mul_re_out(441),
            data_re_in(26) => mul_re_out(442),
            data_re_in(27) => mul_re_out(443),
            data_re_in(28) => mul_re_out(444),
            data_re_in(29) => mul_re_out(445),
            data_re_in(30) => mul_re_out(446),
            data_re_in(31) => mul_re_out(447),
            data_im_in(0) => mul_im_out(416),
            data_im_in(1) => mul_im_out(417),
            data_im_in(2) => mul_im_out(418),
            data_im_in(3) => mul_im_out(419),
            data_im_in(4) => mul_im_out(420),
            data_im_in(5) => mul_im_out(421),
            data_im_in(6) => mul_im_out(422),
            data_im_in(7) => mul_im_out(423),
            data_im_in(8) => mul_im_out(424),
            data_im_in(9) => mul_im_out(425),
            data_im_in(10) => mul_im_out(426),
            data_im_in(11) => mul_im_out(427),
            data_im_in(12) => mul_im_out(428),
            data_im_in(13) => mul_im_out(429),
            data_im_in(14) => mul_im_out(430),
            data_im_in(15) => mul_im_out(431),
            data_im_in(16) => mul_im_out(432),
            data_im_in(17) => mul_im_out(433),
            data_im_in(18) => mul_im_out(434),
            data_im_in(19) => mul_im_out(435),
            data_im_in(20) => mul_im_out(436),
            data_im_in(21) => mul_im_out(437),
            data_im_in(22) => mul_im_out(438),
            data_im_in(23) => mul_im_out(439),
            data_im_in(24) => mul_im_out(440),
            data_im_in(25) => mul_im_out(441),
            data_im_in(26) => mul_im_out(442),
            data_im_in(27) => mul_im_out(443),
            data_im_in(28) => mul_im_out(444),
            data_im_in(29) => mul_im_out(445),
            data_im_in(30) => mul_im_out(446),
            data_im_in(31) => mul_im_out(447),
            data_re_out(0) => data_re_out(13),
            data_re_out(1) => data_re_out(29),
            data_re_out(2) => data_re_out(45),
            data_re_out(3) => data_re_out(61),
            data_re_out(4) => data_re_out(77),
            data_re_out(5) => data_re_out(93),
            data_re_out(6) => data_re_out(109),
            data_re_out(7) => data_re_out(125),
            data_re_out(8) => data_re_out(141),
            data_re_out(9) => data_re_out(157),
            data_re_out(10) => data_re_out(173),
            data_re_out(11) => data_re_out(189),
            data_re_out(12) => data_re_out(205),
            data_re_out(13) => data_re_out(221),
            data_re_out(14) => data_re_out(237),
            data_re_out(15) => data_re_out(253),
            data_re_out(16) => data_re_out(269),
            data_re_out(17) => data_re_out(285),
            data_re_out(18) => data_re_out(301),
            data_re_out(19) => data_re_out(317),
            data_re_out(20) => data_re_out(333),
            data_re_out(21) => data_re_out(349),
            data_re_out(22) => data_re_out(365),
            data_re_out(23) => data_re_out(381),
            data_re_out(24) => data_re_out(397),
            data_re_out(25) => data_re_out(413),
            data_re_out(26) => data_re_out(429),
            data_re_out(27) => data_re_out(445),
            data_re_out(28) => data_re_out(461),
            data_re_out(29) => data_re_out(477),
            data_re_out(30) => data_re_out(493),
            data_re_out(31) => data_re_out(509),
            data_im_out(0) => data_im_out(13),
            data_im_out(1) => data_im_out(29),
            data_im_out(2) => data_im_out(45),
            data_im_out(3) => data_im_out(61),
            data_im_out(4) => data_im_out(77),
            data_im_out(5) => data_im_out(93),
            data_im_out(6) => data_im_out(109),
            data_im_out(7) => data_im_out(125),
            data_im_out(8) => data_im_out(141),
            data_im_out(9) => data_im_out(157),
            data_im_out(10) => data_im_out(173),
            data_im_out(11) => data_im_out(189),
            data_im_out(12) => data_im_out(205),
            data_im_out(13) => data_im_out(221),
            data_im_out(14) => data_im_out(237),
            data_im_out(15) => data_im_out(253),
            data_im_out(16) => data_im_out(269),
            data_im_out(17) => data_im_out(285),
            data_im_out(18) => data_im_out(301),
            data_im_out(19) => data_im_out(317),
            data_im_out(20) => data_im_out(333),
            data_im_out(21) => data_im_out(349),
            data_im_out(22) => data_im_out(365),
            data_im_out(23) => data_im_out(381),
            data_im_out(24) => data_im_out(397),
            data_im_out(25) => data_im_out(413),
            data_im_out(26) => data_im_out(429),
            data_im_out(27) => data_im_out(445),
            data_im_out(28) => data_im_out(461),
            data_im_out(29) => data_im_out(477),
            data_im_out(30) => data_im_out(493),
            data_im_out(31) => data_im_out(509)
        );           

    URFFT_PT32_14 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(448),
            data_re_in(1) => mul_re_out(449),
            data_re_in(2) => mul_re_out(450),
            data_re_in(3) => mul_re_out(451),
            data_re_in(4) => mul_re_out(452),
            data_re_in(5) => mul_re_out(453),
            data_re_in(6) => mul_re_out(454),
            data_re_in(7) => mul_re_out(455),
            data_re_in(8) => mul_re_out(456),
            data_re_in(9) => mul_re_out(457),
            data_re_in(10) => mul_re_out(458),
            data_re_in(11) => mul_re_out(459),
            data_re_in(12) => mul_re_out(460),
            data_re_in(13) => mul_re_out(461),
            data_re_in(14) => mul_re_out(462),
            data_re_in(15) => mul_re_out(463),
            data_re_in(16) => mul_re_out(464),
            data_re_in(17) => mul_re_out(465),
            data_re_in(18) => mul_re_out(466),
            data_re_in(19) => mul_re_out(467),
            data_re_in(20) => mul_re_out(468),
            data_re_in(21) => mul_re_out(469),
            data_re_in(22) => mul_re_out(470),
            data_re_in(23) => mul_re_out(471),
            data_re_in(24) => mul_re_out(472),
            data_re_in(25) => mul_re_out(473),
            data_re_in(26) => mul_re_out(474),
            data_re_in(27) => mul_re_out(475),
            data_re_in(28) => mul_re_out(476),
            data_re_in(29) => mul_re_out(477),
            data_re_in(30) => mul_re_out(478),
            data_re_in(31) => mul_re_out(479),
            data_im_in(0) => mul_im_out(448),
            data_im_in(1) => mul_im_out(449),
            data_im_in(2) => mul_im_out(450),
            data_im_in(3) => mul_im_out(451),
            data_im_in(4) => mul_im_out(452),
            data_im_in(5) => mul_im_out(453),
            data_im_in(6) => mul_im_out(454),
            data_im_in(7) => mul_im_out(455),
            data_im_in(8) => mul_im_out(456),
            data_im_in(9) => mul_im_out(457),
            data_im_in(10) => mul_im_out(458),
            data_im_in(11) => mul_im_out(459),
            data_im_in(12) => mul_im_out(460),
            data_im_in(13) => mul_im_out(461),
            data_im_in(14) => mul_im_out(462),
            data_im_in(15) => mul_im_out(463),
            data_im_in(16) => mul_im_out(464),
            data_im_in(17) => mul_im_out(465),
            data_im_in(18) => mul_im_out(466),
            data_im_in(19) => mul_im_out(467),
            data_im_in(20) => mul_im_out(468),
            data_im_in(21) => mul_im_out(469),
            data_im_in(22) => mul_im_out(470),
            data_im_in(23) => mul_im_out(471),
            data_im_in(24) => mul_im_out(472),
            data_im_in(25) => mul_im_out(473),
            data_im_in(26) => mul_im_out(474),
            data_im_in(27) => mul_im_out(475),
            data_im_in(28) => mul_im_out(476),
            data_im_in(29) => mul_im_out(477),
            data_im_in(30) => mul_im_out(478),
            data_im_in(31) => mul_im_out(479),
            data_re_out(0) => data_re_out(14),
            data_re_out(1) => data_re_out(30),
            data_re_out(2) => data_re_out(46),
            data_re_out(3) => data_re_out(62),
            data_re_out(4) => data_re_out(78),
            data_re_out(5) => data_re_out(94),
            data_re_out(6) => data_re_out(110),
            data_re_out(7) => data_re_out(126),
            data_re_out(8) => data_re_out(142),
            data_re_out(9) => data_re_out(158),
            data_re_out(10) => data_re_out(174),
            data_re_out(11) => data_re_out(190),
            data_re_out(12) => data_re_out(206),
            data_re_out(13) => data_re_out(222),
            data_re_out(14) => data_re_out(238),
            data_re_out(15) => data_re_out(254),
            data_re_out(16) => data_re_out(270),
            data_re_out(17) => data_re_out(286),
            data_re_out(18) => data_re_out(302),
            data_re_out(19) => data_re_out(318),
            data_re_out(20) => data_re_out(334),
            data_re_out(21) => data_re_out(350),
            data_re_out(22) => data_re_out(366),
            data_re_out(23) => data_re_out(382),
            data_re_out(24) => data_re_out(398),
            data_re_out(25) => data_re_out(414),
            data_re_out(26) => data_re_out(430),
            data_re_out(27) => data_re_out(446),
            data_re_out(28) => data_re_out(462),
            data_re_out(29) => data_re_out(478),
            data_re_out(30) => data_re_out(494),
            data_re_out(31) => data_re_out(510),
            data_im_out(0) => data_im_out(14),
            data_im_out(1) => data_im_out(30),
            data_im_out(2) => data_im_out(46),
            data_im_out(3) => data_im_out(62),
            data_im_out(4) => data_im_out(78),
            data_im_out(5) => data_im_out(94),
            data_im_out(6) => data_im_out(110),
            data_im_out(7) => data_im_out(126),
            data_im_out(8) => data_im_out(142),
            data_im_out(9) => data_im_out(158),
            data_im_out(10) => data_im_out(174),
            data_im_out(11) => data_im_out(190),
            data_im_out(12) => data_im_out(206),
            data_im_out(13) => data_im_out(222),
            data_im_out(14) => data_im_out(238),
            data_im_out(15) => data_im_out(254),
            data_im_out(16) => data_im_out(270),
            data_im_out(17) => data_im_out(286),
            data_im_out(18) => data_im_out(302),
            data_im_out(19) => data_im_out(318),
            data_im_out(20) => data_im_out(334),
            data_im_out(21) => data_im_out(350),
            data_im_out(22) => data_im_out(366),
            data_im_out(23) => data_im_out(382),
            data_im_out(24) => data_im_out(398),
            data_im_out(25) => data_im_out(414),
            data_im_out(26) => data_im_out(430),
            data_im_out(27) => data_im_out(446),
            data_im_out(28) => data_im_out(462),
            data_im_out(29) => data_im_out(478),
            data_im_out(30) => data_im_out(494),
            data_im_out(31) => data_im_out(510)
        );           

    URFFT_PT32_15 : fft_pt32
    generic map(
        ctrl_start => (ctrl_start+4) mod 16
    )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(4 DOWNTO 0),
            ctrl_delay => ctrl_delay,
            data_re_in(0) => mul_re_out(480),
            data_re_in(1) => mul_re_out(481),
            data_re_in(2) => mul_re_out(482),
            data_re_in(3) => mul_re_out(483),
            data_re_in(4) => mul_re_out(484),
            data_re_in(5) => mul_re_out(485),
            data_re_in(6) => mul_re_out(486),
            data_re_in(7) => mul_re_out(487),
            data_re_in(8) => mul_re_out(488),
            data_re_in(9) => mul_re_out(489),
            data_re_in(10) => mul_re_out(490),
            data_re_in(11) => mul_re_out(491),
            data_re_in(12) => mul_re_out(492),
            data_re_in(13) => mul_re_out(493),
            data_re_in(14) => mul_re_out(494),
            data_re_in(15) => mul_re_out(495),
            data_re_in(16) => mul_re_out(496),
            data_re_in(17) => mul_re_out(497),
            data_re_in(18) => mul_re_out(498),
            data_re_in(19) => mul_re_out(499),
            data_re_in(20) => mul_re_out(500),
            data_re_in(21) => mul_re_out(501),
            data_re_in(22) => mul_re_out(502),
            data_re_in(23) => mul_re_out(503),
            data_re_in(24) => mul_re_out(504),
            data_re_in(25) => mul_re_out(505),
            data_re_in(26) => mul_re_out(506),
            data_re_in(27) => mul_re_out(507),
            data_re_in(28) => mul_re_out(508),
            data_re_in(29) => mul_re_out(509),
            data_re_in(30) => mul_re_out(510),
            data_re_in(31) => mul_re_out(511),
            data_im_in(0) => mul_im_out(480),
            data_im_in(1) => mul_im_out(481),
            data_im_in(2) => mul_im_out(482),
            data_im_in(3) => mul_im_out(483),
            data_im_in(4) => mul_im_out(484),
            data_im_in(5) => mul_im_out(485),
            data_im_in(6) => mul_im_out(486),
            data_im_in(7) => mul_im_out(487),
            data_im_in(8) => mul_im_out(488),
            data_im_in(9) => mul_im_out(489),
            data_im_in(10) => mul_im_out(490),
            data_im_in(11) => mul_im_out(491),
            data_im_in(12) => mul_im_out(492),
            data_im_in(13) => mul_im_out(493),
            data_im_in(14) => mul_im_out(494),
            data_im_in(15) => mul_im_out(495),
            data_im_in(16) => mul_im_out(496),
            data_im_in(17) => mul_im_out(497),
            data_im_in(18) => mul_im_out(498),
            data_im_in(19) => mul_im_out(499),
            data_im_in(20) => mul_im_out(500),
            data_im_in(21) => mul_im_out(501),
            data_im_in(22) => mul_im_out(502),
            data_im_in(23) => mul_im_out(503),
            data_im_in(24) => mul_im_out(504),
            data_im_in(25) => mul_im_out(505),
            data_im_in(26) => mul_im_out(506),
            data_im_in(27) => mul_im_out(507),
            data_im_in(28) => mul_im_out(508),
            data_im_in(29) => mul_im_out(509),
            data_im_in(30) => mul_im_out(510),
            data_im_in(31) => mul_im_out(511),
            data_re_out(0) => data_re_out(15),
            data_re_out(1) => data_re_out(31),
            data_re_out(2) => data_re_out(47),
            data_re_out(3) => data_re_out(63),
            data_re_out(4) => data_re_out(79),
            data_re_out(5) => data_re_out(95),
            data_re_out(6) => data_re_out(111),
            data_re_out(7) => data_re_out(127),
            data_re_out(8) => data_re_out(143),
            data_re_out(9) => data_re_out(159),
            data_re_out(10) => data_re_out(175),
            data_re_out(11) => data_re_out(191),
            data_re_out(12) => data_re_out(207),
            data_re_out(13) => data_re_out(223),
            data_re_out(14) => data_re_out(239),
            data_re_out(15) => data_re_out(255),
            data_re_out(16) => data_re_out(271),
            data_re_out(17) => data_re_out(287),
            data_re_out(18) => data_re_out(303),
            data_re_out(19) => data_re_out(319),
            data_re_out(20) => data_re_out(335),
            data_re_out(21) => data_re_out(351),
            data_re_out(22) => data_re_out(367),
            data_re_out(23) => data_re_out(383),
            data_re_out(24) => data_re_out(399),
            data_re_out(25) => data_re_out(415),
            data_re_out(26) => data_re_out(431),
            data_re_out(27) => data_re_out(447),
            data_re_out(28) => data_re_out(463),
            data_re_out(29) => data_re_out(479),
            data_re_out(30) => data_re_out(495),
            data_re_out(31) => data_re_out(511),
            data_im_out(0) => data_im_out(15),
            data_im_out(1) => data_im_out(31),
            data_im_out(2) => data_im_out(47),
            data_im_out(3) => data_im_out(63),
            data_im_out(4) => data_im_out(79),
            data_im_out(5) => data_im_out(95),
            data_im_out(6) => data_im_out(111),
            data_im_out(7) => data_im_out(127),
            data_im_out(8) => data_im_out(143),
            data_im_out(9) => data_im_out(159),
            data_im_out(10) => data_im_out(175),
            data_im_out(11) => data_im_out(191),
            data_im_out(12) => data_im_out(207),
            data_im_out(13) => data_im_out(223),
            data_im_out(14) => data_im_out(239),
            data_im_out(15) => data_im_out(255),
            data_im_out(16) => data_im_out(271),
            data_im_out(17) => data_im_out(287),
            data_im_out(18) => data_im_out(303),
            data_im_out(19) => data_im_out(319),
            data_im_out(20) => data_im_out(335),
            data_im_out(21) => data_im_out(351),
            data_im_out(22) => data_im_out(367),
            data_im_out(23) => data_im_out(383),
            data_im_out(24) => data_im_out(399),
            data_im_out(25) => data_im_out(415),
            data_im_out(26) => data_im_out(431),
            data_im_out(27) => data_im_out(447),
            data_im_out(28) => data_im_out(463),
            data_im_out(29) => data_im_out(479),
            data_im_out(30) => data_im_out(495),
            data_im_out(31) => data_im_out(511)
        );           


    --- multipliers
 
    UMUL_0 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(0),
            data_im_in => first_stage_im_out(0),
            data_re_out => mul_re_out(0),
            data_im_out => mul_im_out(0)
        );

 
    UMUL_1 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(1),
            data_im_in => first_stage_im_out(1),
            data_re_out => mul_re_out(1),
            data_im_out => mul_im_out(1)
        );

 
    UMUL_2 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(2),
            data_im_in => first_stage_im_out(2),
            data_re_out => mul_re_out(2),
            data_im_out => mul_im_out(2)
        );

 
    UMUL_3 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(3),
            data_im_in => first_stage_im_out(3),
            data_re_out => mul_re_out(3),
            data_im_out => mul_im_out(3)
        );

 
    UMUL_4 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(4),
            data_im_in => first_stage_im_out(4),
            data_re_out => mul_re_out(4),
            data_im_out => mul_im_out(4)
        );

 
    UMUL_5 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(5),
            data_im_in => first_stage_im_out(5),
            data_re_out => mul_re_out(5),
            data_im_out => mul_im_out(5)
        );

 
    UMUL_6 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(6),
            data_im_in => first_stage_im_out(6),
            data_re_out => mul_re_out(6),
            data_im_out => mul_im_out(6)
        );

 
    UMUL_7 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(7),
            data_im_in => first_stage_im_out(7),
            data_re_out => mul_re_out(7),
            data_im_out => mul_im_out(7)
        );

 
    UMUL_8 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(8),
            data_im_in => first_stage_im_out(8),
            data_re_out => mul_re_out(8),
            data_im_out => mul_im_out(8)
        );

 
    UMUL_9 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(9),
            data_im_in => first_stage_im_out(9),
            data_re_out => mul_re_out(9),
            data_im_out => mul_im_out(9)
        );

 
    UMUL_10 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(10),
            data_im_in => first_stage_im_out(10),
            data_re_out => mul_re_out(10),
            data_im_out => mul_im_out(10)
        );

 
    UMUL_11 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(11),
            data_im_in => first_stage_im_out(11),
            data_re_out => mul_re_out(11),
            data_im_out => mul_im_out(11)
        );

 
    UMUL_12 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(12),
            data_im_in => first_stage_im_out(12),
            data_re_out => mul_re_out(12),
            data_im_out => mul_im_out(12)
        );

 
    UMUL_13 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(13),
            data_im_in => first_stage_im_out(13),
            data_re_out => mul_re_out(13),
            data_im_out => mul_im_out(13)
        );

 
    UMUL_14 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(14),
            data_im_in => first_stage_im_out(14),
            data_re_out => mul_re_out(14),
            data_im_out => mul_im_out(14)
        );

 
    UMUL_15 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(15),
            data_im_in => first_stage_im_out(15),
            data_re_out => mul_re_out(15),
            data_im_out => mul_im_out(15)
        );

 
    UMUL_16 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(16),
            data_im_in => first_stage_im_out(16),
            data_re_out => mul_re_out(16),
            data_im_out => mul_im_out(16)
        );

 
    UMUL_17 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(17),
            data_im_in => first_stage_im_out(17),
            data_re_out => mul_re_out(17),
            data_im_out => mul_im_out(17)
        );

 
    UMUL_18 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(18),
            data_im_in => first_stage_im_out(18),
            data_re_out => mul_re_out(18),
            data_im_out => mul_im_out(18)
        );

 
    UMUL_19 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(19),
            data_im_in => first_stage_im_out(19),
            data_re_out => mul_re_out(19),
            data_im_out => mul_im_out(19)
        );

 
    UMUL_20 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(20),
            data_im_in => first_stage_im_out(20),
            data_re_out => mul_re_out(20),
            data_im_out => mul_im_out(20)
        );

 
    UMUL_21 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(21),
            data_im_in => first_stage_im_out(21),
            data_re_out => mul_re_out(21),
            data_im_out => mul_im_out(21)
        );

 
    UMUL_22 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(22),
            data_im_in => first_stage_im_out(22),
            data_re_out => mul_re_out(22),
            data_im_out => mul_im_out(22)
        );

 
    UMUL_23 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(23),
            data_im_in => first_stage_im_out(23),
            data_re_out => mul_re_out(23),
            data_im_out => mul_im_out(23)
        );

 
    UMUL_24 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(24),
            data_im_in => first_stage_im_out(24),
            data_re_out => mul_re_out(24),
            data_im_out => mul_im_out(24)
        );

 
    UMUL_25 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(25),
            data_im_in => first_stage_im_out(25),
            data_re_out => mul_re_out(25),
            data_im_out => mul_im_out(25)
        );

 
    UMUL_26 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(26),
            data_im_in => first_stage_im_out(26),
            data_re_out => mul_re_out(26),
            data_im_out => mul_im_out(26)
        );

 
    UMUL_27 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(27),
            data_im_in => first_stage_im_out(27),
            data_re_out => mul_re_out(27),
            data_im_out => mul_im_out(27)
        );

 
    UMUL_28 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(28),
            data_im_in => first_stage_im_out(28),
            data_re_out => mul_re_out(28),
            data_im_out => mul_im_out(28)
        );

 
    UMUL_29 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(29),
            data_im_in => first_stage_im_out(29),
            data_re_out => mul_re_out(29),
            data_im_out => mul_im_out(29)
        );

 
    UMUL_30 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(30),
            data_im_in => first_stage_im_out(30),
            data_re_out => mul_re_out(30),
            data_im_out => mul_im_out(30)
        );

 
    UMUL_31 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(31),
            data_im_in => first_stage_im_out(31),
            data_re_out => mul_re_out(31),
            data_im_out => mul_im_out(31)
        );

 
    UMUL_32 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(32),
            data_im_in => first_stage_im_out(32),
            data_re_out => mul_re_out(32),
            data_im_out => mul_im_out(32)
        );

 
    UMUL_33 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(33),
            data_im_in => first_stage_im_out(33),
            re_multiplicator => "0011111111111111", --- 0.999938964844 + j-0.0122680664062
            im_multiplicator => "1111111100110111",
            data_re_out => mul_re_out(33),
            data_im_out => mul_im_out(33)
        );

 
    UMUL_34 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(34),
            data_im_in => first_stage_im_out(34),
            re_multiplicator => "0011111111111011", --- 0.999694824219 + j-0.0245361328125
            im_multiplicator => "1111111001101110",
            data_re_out => mul_re_out(34),
            data_im_out => mul_im_out(34)
        );

 
    UMUL_35 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(35),
            data_im_in => first_stage_im_out(35),
            re_multiplicator => "0011111111110101", --- 0.999328613281 + j-0.0368041992188
            im_multiplicator => "1111110110100101",
            data_re_out => mul_re_out(35),
            data_im_out => mul_im_out(35)
        );

 
    UMUL_36 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(36),
            data_im_in => first_stage_im_out(36),
            re_multiplicator => "0011111111101100", --- 0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(36),
            data_im_out => mul_im_out(36)
        );

 
    UMUL_37 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(37),
            data_im_in => first_stage_im_out(37),
            re_multiplicator => "0011111111100001", --- 0.998107910156 + j-0.0613403320312
            im_multiplicator => "1111110000010011",
            data_re_out => mul_re_out(37),
            data_im_out => mul_im_out(37)
        );

 
    UMUL_38 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(38),
            data_im_in => first_stage_im_out(38),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(38),
            data_im_out => mul_im_out(38)
        );

 
    UMUL_39 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(39),
            data_im_in => first_stage_im_out(39),
            re_multiplicator => "0011111111000100", --- 0.996337890625 + j-0.0858154296875
            im_multiplicator => "1111101010000010",
            data_re_out => mul_re_out(39),
            data_im_out => mul_im_out(39)
        );

 
    UMUL_40 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(40),
            data_im_in => first_stage_im_out(40),
            re_multiplicator => "0011111110110001", --- 0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(40),
            data_im_out => mul_im_out(40)
        );

 
    UMUL_41 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(41),
            data_im_in => first_stage_im_out(41),
            re_multiplicator => "0011111110011100", --- 0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(41),
            data_im_out => mul_im_out(41)
        );

 
    UMUL_42 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(42),
            data_im_in => first_stage_im_out(42),
            re_multiplicator => "0011111110000101", --- 0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(42),
            data_im_out => mul_im_out(42)
        );

 
    UMUL_43 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(43),
            data_im_in => first_stage_im_out(43),
            re_multiplicator => "0011111101101011", --- 0.990905761719 + j-0.134582519531
            im_multiplicator => "1111011101100011",
            data_re_out => mul_re_out(43),
            data_im_out => mul_im_out(43)
        );

 
    UMUL_44 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(44),
            data_im_in => first_stage_im_out(44),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(44),
            data_im_out => mul_im_out(44)
        );

 
    UMUL_45 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(45),
            data_im_in => first_stage_im_out(45),
            re_multiplicator => "0011111100110000", --- 0.9873046875 + j-0.158874511719
            im_multiplicator => "1111010111010101",
            data_re_out => mul_re_out(45),
            data_im_out => mul_im_out(45)
        );

 
    UMUL_46 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(46),
            data_im_in => first_stage_im_out(46),
            re_multiplicator => "0011111100001111", --- 0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(46),
            data_im_out => mul_im_out(46)
        );

 
    UMUL_47 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(47),
            data_im_in => first_stage_im_out(47),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(47),
            data_im_out => mul_im_out(47)
        );

 
    UMUL_48 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(48),
            data_im_in => first_stage_im_out(48),
            re_multiplicator => "0011111011000101", --- 0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(48),
            data_im_out => mul_im_out(48)
        );

 
    UMUL_49 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(49),
            data_im_in => first_stage_im_out(49),
            re_multiplicator => "0011111010011101", --- 0.978332519531 + j-0.207092285156
            im_multiplicator => "1111001010111111",
            data_re_out => mul_re_out(49),
            data_im_out => mul_im_out(49)
        );

 
    UMUL_50 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(50),
            data_im_in => first_stage_im_out(50),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(50),
            data_im_out => mul_im_out(50)
        );

 
    UMUL_51 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(51),
            data_im_in => first_stage_im_out(51),
            re_multiplicator => "0011111001000101", --- 0.972961425781 + j-0.231079101562
            im_multiplicator => "1111000100110110",
            data_re_out => mul_re_out(51),
            data_im_out => mul_im_out(51)
        );

 
    UMUL_52 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(52),
            data_im_in => first_stage_im_out(52),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(52),
            data_im_out => mul_im_out(52)
        );

 
    UMUL_53 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(53),
            data_im_in => first_stage_im_out(53),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(53),
            data_im_out => mul_im_out(53)
        );

 
    UMUL_54 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(54),
            data_im_in => first_stage_im_out(54),
            re_multiplicator => "0011110110101111", --- 0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(54),
            data_im_out => mul_im_out(54)
        );

 
    UMUL_55 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(55),
            data_im_in => first_stage_im_out(55),
            re_multiplicator => "0011110101111000", --- 0.96044921875 + j-0.278503417969
            im_multiplicator => "1110111000101101",
            data_re_out => mul_re_out(55),
            data_im_out => mul_im_out(55)
        );

 
    UMUL_56 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(56),
            data_im_in => first_stage_im_out(56),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(56),
            data_im_out => mul_im_out(56)
        );

 
    UMUL_57 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(57),
            data_im_in => first_stage_im_out(57),
            re_multiplicator => "0011110100000011", --- 0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(57),
            data_im_out => mul_im_out(57)
        );

 
    UMUL_58 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(58),
            data_im_in => first_stage_im_out(58),
            re_multiplicator => "0011110011000101", --- 0.949523925781 + j-0.313659667969
            im_multiplicator => "1110101111101101",
            data_re_out => mul_re_out(58),
            data_im_out => mul_im_out(58)
        );

 
    UMUL_59 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(59),
            data_im_in => first_stage_im_out(59),
            re_multiplicator => "0011110010000101", --- 0.945617675781 + j-0.325317382812
            im_multiplicator => "1110101100101110",
            data_re_out => mul_re_out(59),
            data_im_out => mul_im_out(59)
        );

 
    UMUL_60 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(60),
            data_im_in => first_stage_im_out(60),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(60),
            data_im_out => mul_im_out(60)
        );

 
    UMUL_61 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(61),
            data_im_in => first_stage_im_out(61),
            re_multiplicator => "0011101111111101", --- 0.937316894531 + j-0.348388671875
            im_multiplicator => "1110100110110100",
            data_re_out => mul_re_out(61),
            data_im_out => mul_im_out(61)
        );

 
    UMUL_62 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(62),
            data_im_in => first_stage_im_out(62),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(62),
            data_im_out => mul_im_out(62)
        );

 
    UMUL_63 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(63),
            data_im_in => first_stage_im_out(63),
            re_multiplicator => "0011101101101101", --- 0.928527832031 + j-0.371337890625
            im_multiplicator => "1110100000111100",
            data_re_out => mul_re_out(63),
            data_im_out => mul_im_out(63)
        );

 
    UMUL_64 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(64),
            data_im_in => first_stage_im_out(64),
            data_re_out => mul_re_out(64),
            data_im_out => mul_im_out(64)
        );

 
    UMUL_65 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(65),
            data_im_in => first_stage_im_out(65),
            re_multiplicator => "0011111111111011", --- 0.999694824219 + j-0.0245361328125
            im_multiplicator => "1111111001101110",
            data_re_out => mul_re_out(65),
            data_im_out => mul_im_out(65)
        );

 
    UMUL_66 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(66),
            data_im_in => first_stage_im_out(66),
            re_multiplicator => "0011111111101100", --- 0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(66),
            data_im_out => mul_im_out(66)
        );

 
    UMUL_67 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(67),
            data_im_in => first_stage_im_out(67),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(67),
            data_im_out => mul_im_out(67)
        );

 
    UMUL_68 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(68),
            data_im_in => first_stage_im_out(68),
            re_multiplicator => "0011111110110001", --- 0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(68),
            data_im_out => mul_im_out(68)
        );

 
    UMUL_69 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(69),
            data_im_in => first_stage_im_out(69),
            re_multiplicator => "0011111110000101", --- 0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(69),
            data_im_out => mul_im_out(69)
        );

 
    UMUL_70 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(70),
            data_im_in => first_stage_im_out(70),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(70),
            data_im_out => mul_im_out(70)
        );

 
    UMUL_71 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(71),
            data_im_in => first_stage_im_out(71),
            re_multiplicator => "0011111100001111", --- 0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(71),
            data_im_out => mul_im_out(71)
        );

 
    UMUL_72 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(72),
            data_im_in => first_stage_im_out(72),
            re_multiplicator => "0011111011000101", --- 0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(72),
            data_im_out => mul_im_out(72)
        );

 
    UMUL_73 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(73),
            data_im_in => first_stage_im_out(73),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(73),
            data_im_out => mul_im_out(73)
        );

 
    UMUL_74 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(74),
            data_im_in => first_stage_im_out(74),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(74),
            data_im_out => mul_im_out(74)
        );

 
    UMUL_75 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(75),
            data_im_in => first_stage_im_out(75),
            re_multiplicator => "0011110110101111", --- 0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(75),
            data_im_out => mul_im_out(75)
        );

 
    UMUL_76 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(76),
            data_im_in => first_stage_im_out(76),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(76),
            data_im_out => mul_im_out(76)
        );

 
    UMUL_77 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(77),
            data_im_in => first_stage_im_out(77),
            re_multiplicator => "0011110011000101", --- 0.949523925781 + j-0.313659667969
            im_multiplicator => "1110101111101101",
            data_re_out => mul_re_out(77),
            data_im_out => mul_im_out(77)
        );

 
    UMUL_78 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(78),
            data_im_in => first_stage_im_out(78),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(78),
            data_im_out => mul_im_out(78)
        );

 
    UMUL_79 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(79),
            data_im_in => first_stage_im_out(79),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(79),
            data_im_out => mul_im_out(79)
        );

 
    UMUL_80 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(80),
            data_im_in => first_stage_im_out(80),
            re_multiplicator => "0011101100100001", --- 0.923889160156 + j-0.382690429688
            im_multiplicator => "1110011110000010",
            data_re_out => mul_re_out(80),
            data_im_out => mul_im_out(80)
        );

 
    UMUL_81 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(81),
            data_im_in => first_stage_im_out(81),
            re_multiplicator => "0011101010000010", --- 0.914184570312 + j-0.405212402344
            im_multiplicator => "1110011000010001",
            data_re_out => mul_re_out(81),
            data_im_out => mul_im_out(81)
        );

 
    UMUL_82 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(82),
            data_im_in => first_stage_im_out(82),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(82),
            data_im_out => mul_im_out(82)
        );

 
    UMUL_83 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(83),
            data_im_in => first_stage_im_out(83),
            re_multiplicator => "0011100100101011", --- 0.893249511719 + j-0.449584960938
            im_multiplicator => "1110001100111010",
            data_re_out => mul_re_out(83),
            data_im_out => mul_im_out(83)
        );

 
    UMUL_84 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(84),
            data_im_in => first_stage_im_out(84),
            re_multiplicator => "0011100001110001", --- 0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(84),
            data_im_out => mul_im_out(84)
        );

 
    UMUL_85 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(85),
            data_im_in => first_stage_im_out(85),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(85),
            data_im_out => mul_im_out(85)
        );

 
    UMUL_86 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(86),
            data_im_in => first_stage_im_out(86),
            re_multiplicator => "0011011011100101", --- 0.857727050781 + j-0.514099121094
            im_multiplicator => "1101111100011001",
            data_re_out => mul_re_out(86),
            data_im_out => mul_im_out(86)
        );

 
    UMUL_87 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(87),
            data_im_in => first_stage_im_out(87),
            re_multiplicator => "0011011000010010", --- 0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(87),
            data_im_out => mul_im_out(87)
        );

 
    UMUL_88 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(88),
            data_im_in => first_stage_im_out(88),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(88),
            data_im_out => mul_im_out(88)
        );

 
    UMUL_89 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(89),
            data_im_in => first_stage_im_out(89),
            re_multiplicator => "0011010001010011", --- 0.817565917969 + j-0.575805664062
            im_multiplicator => "1101101100100110",
            data_re_out => mul_re_out(89),
            data_im_out => mul_im_out(89)
        );

 
    UMUL_90 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(90),
            data_im_in => first_stage_im_out(90),
            re_multiplicator => "0011001101101000", --- 0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(90),
            data_im_out => mul_im_out(90)
        );

 
    UMUL_91 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(91),
            data_im_in => first_stage_im_out(91),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(91),
            data_im_out => mul_im_out(91)
        );

 
    UMUL_92 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(92),
            data_im_in => first_stage_im_out(92),
            re_multiplicator => "0011000101111001", --- 0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(92),
            data_im_out => mul_im_out(92)
        );

 
    UMUL_93 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(93),
            data_im_in => first_stage_im_out(93),
            re_multiplicator => "0011000001110110", --- 0.757202148438 + j-0.653198242188
            im_multiplicator => "1101011000110010",
            data_re_out => mul_re_out(93),
            data_im_out => mul_im_out(93)
        );

 
    UMUL_94 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(94),
            data_im_in => first_stage_im_out(94),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(94),
            data_im_out => mul_im_out(94)
        );

 
    UMUL_95 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(95),
            data_im_in => first_stage_im_out(95),
            re_multiplicator => "0010111001011010", --- 0.724243164062 + j-0.689514160156
            im_multiplicator => "1101001111011111",
            data_re_out => mul_re_out(95),
            data_im_out => mul_im_out(95)
        );

 
    UMUL_96 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(96),
            data_im_in => first_stage_im_out(96),
            data_re_out => mul_re_out(96),
            data_im_out => mul_im_out(96)
        );

 
    UMUL_97 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(97),
            data_im_in => first_stage_im_out(97),
            re_multiplicator => "0011111111110101", --- 0.999328613281 + j-0.0368041992188
            im_multiplicator => "1111110110100101",
            data_re_out => mul_re_out(97),
            data_im_out => mul_im_out(97)
        );

 
    UMUL_98 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(98),
            data_im_in => first_stage_im_out(98),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(98),
            data_im_out => mul_im_out(98)
        );

 
    UMUL_99 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(99),
            data_im_in => first_stage_im_out(99),
            re_multiplicator => "0011111110011100", --- 0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(99),
            data_im_out => mul_im_out(99)
        );

 
    UMUL_100 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(100),
            data_im_in => first_stage_im_out(100),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(100),
            data_im_out => mul_im_out(100)
        );

 
    UMUL_101 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(101),
            data_im_in => first_stage_im_out(101),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(101),
            data_im_out => mul_im_out(101)
        );

 
    UMUL_102 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(102),
            data_im_in => first_stage_im_out(102),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(102),
            data_im_out => mul_im_out(102)
        );

 
    UMUL_103 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(103),
            data_im_in => first_stage_im_out(103),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(103),
            data_im_out => mul_im_out(103)
        );

 
    UMUL_104 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(104),
            data_im_in => first_stage_im_out(104),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(104),
            data_im_out => mul_im_out(104)
        );

 
    UMUL_105 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(105),
            data_im_in => first_stage_im_out(105),
            re_multiplicator => "0011110010000101", --- 0.945617675781 + j-0.325317382812
            im_multiplicator => "1110101100101110",
            data_re_out => mul_re_out(105),
            data_im_out => mul_im_out(105)
        );

 
    UMUL_106 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(106),
            data_im_in => first_stage_im_out(106),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(106),
            data_im_out => mul_im_out(106)
        );

 
    UMUL_107 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(107),
            data_im_in => first_stage_im_out(107),
            re_multiplicator => "0011101011010011", --- 0.919128417969 + j-0.393981933594
            im_multiplicator => "1110011011001001",
            data_re_out => mul_re_out(107),
            data_im_out => mul_im_out(107)
        );

 
    UMUL_108 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(108),
            data_im_in => first_stage_im_out(108),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(108),
            data_im_out => mul_im_out(108)
        );

 
    UMUL_109 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(109),
            data_im_in => first_stage_im_out(109),
            re_multiplicator => "0011100011001111", --- 0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(109),
            data_im_out => mul_im_out(109)
        );

 
    UMUL_110 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(110),
            data_im_in => first_stage_im_out(110),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(110),
            data_im_out => mul_im_out(110)
        );

 
    UMUL_111 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(111),
            data_im_in => first_stage_im_out(111),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(111),
            data_im_out => mul_im_out(111)
        );

 
    UMUL_112 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(112),
            data_im_in => first_stage_im_out(112),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(112),
            data_im_out => mul_im_out(112)
        );

 
    UMUL_113 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(113),
            data_im_in => first_stage_im_out(113),
            re_multiplicator => "0011001111011111", --- 0.810485839844 + j-0.585815429688
            im_multiplicator => "1101101010000010",
            data_re_out => mul_re_out(113),
            data_im_out => mul_im_out(113)
        );

 
    UMUL_114 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(114),
            data_im_in => first_stage_im_out(114),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(114),
            data_im_out => mul_im_out(114)
        );

 
    UMUL_115 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(115),
            data_im_in => first_stage_im_out(115),
            re_multiplicator => "0011000011111001", --- 0.765197753906 + j-0.643859863281
            im_multiplicator => "1101011011001011",
            data_re_out => mul_re_out(115),
            data_im_out => mul_im_out(115)
        );

 
    UMUL_116 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(116),
            data_im_in => first_stage_im_out(116),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(116),
            data_im_out => mul_im_out(116)
        );

 
    UMUL_117 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(117),
            data_im_in => first_stage_im_out(117),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(117),
            data_im_out => mul_im_out(117)
        );

 
    UMUL_118 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(118),
            data_im_in => first_stage_im_out(118),
            re_multiplicator => "0010110000100001", --- 0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(118),
            data_im_out => mul_im_out(118)
        );

 
    UMUL_119 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(119),
            data_im_in => first_stage_im_out(119),
            re_multiplicator => "0010101001100101", --- 0.662414550781 + j-0.749145507812
            im_multiplicator => "1101000000001110",
            data_re_out => mul_re_out(119),
            data_im_out => mul_im_out(119)
        );

 
    UMUL_120 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(120),
            data_im_in => first_stage_im_out(120),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(120),
            data_im_out => mul_im_out(120)
        );

 
    UMUL_121 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(121),
            data_im_in => first_stage_im_out(121),
            re_multiplicator => "0010011011000001", --- 0.605529785156 + j-0.795837402344
            im_multiplicator => "1100110100010001",
            data_re_out => mul_re_out(121),
            data_im_out => mul_im_out(121)
        );

 
    UMUL_122 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(122),
            data_im_in => first_stage_im_out(122),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j-0.817565917969
            im_multiplicator => "1100101110101101",
            data_re_out => mul_re_out(122),
            data_im_out => mul_im_out(122)
        );

 
    UMUL_123 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(123),
            data_im_in => first_stage_im_out(123),
            re_multiplicator => "0010001011100111", --- 0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(123),
            data_im_out => mul_im_out(123)
        );

 
    UMUL_124 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(124),
            data_im_in => first_stage_im_out(124),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(124),
            data_im_out => mul_im_out(124)
        );

 
    UMUL_125 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(125),
            data_im_in => first_stage_im_out(125),
            re_multiplicator => "0001111011011100", --- 0.482177734375 + j-0.876098632812
            im_multiplicator => "1100011111101110",
            data_re_out => mul_re_out(125),
            data_im_out => mul_im_out(125)
        );

 
    UMUL_126 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(126),
            data_im_in => first_stage_im_out(126),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(126),
            data_im_out => mul_im_out(126)
        );

 
    UMUL_127 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(127),
            data_im_in => first_stage_im_out(127),
            re_multiplicator => "0001101010100111", --- 0.416442871094 + j-0.9091796875
            im_multiplicator => "1100010111010000",
            data_re_out => mul_re_out(127),
            data_im_out => mul_im_out(127)
        );

 
    UMUL_128 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(128),
            data_im_in => first_stage_im_out(128),
            data_re_out => mul_re_out(128),
            data_im_out => mul_im_out(128)
        );

 
    UMUL_129 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(129),
            data_im_in => first_stage_im_out(129),
            re_multiplicator => "0011111111101100", --- 0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(129),
            data_im_out => mul_im_out(129)
        );

 
    UMUL_130 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(130),
            data_im_in => first_stage_im_out(130),
            re_multiplicator => "0011111110110001", --- 0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(130),
            data_im_out => mul_im_out(130)
        );

 
    UMUL_131 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(131),
            data_im_in => first_stage_im_out(131),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(131),
            data_im_out => mul_im_out(131)
        );

 
    UMUL_132 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(132),
            data_im_in => first_stage_im_out(132),
            re_multiplicator => "0011111011000101", --- 0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(132),
            data_im_out => mul_im_out(132)
        );

 
    UMUL_133 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(133),
            data_im_in => first_stage_im_out(133),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(133),
            data_im_out => mul_im_out(133)
        );

 
    UMUL_134 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(134),
            data_im_in => first_stage_im_out(134),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(134),
            data_im_out => mul_im_out(134)
        );

 
    UMUL_135 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(135),
            data_im_in => first_stage_im_out(135),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(135),
            data_im_out => mul_im_out(135)
        );

 
    UMUL_136 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(136),
            data_im_in => first_stage_im_out(136),
            re_multiplicator => "0011101100100001", --- 0.923889160156 + j-0.382690429688
            im_multiplicator => "1110011110000010",
            data_re_out => mul_re_out(136),
            data_im_out => mul_im_out(136)
        );

 
    UMUL_137 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(137),
            data_im_in => first_stage_im_out(137),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(137),
            data_im_out => mul_im_out(137)
        );

 
    UMUL_138 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(138),
            data_im_in => first_stage_im_out(138),
            re_multiplicator => "0011100001110001", --- 0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(138),
            data_im_out => mul_im_out(138)
        );

 
    UMUL_139 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(139),
            data_im_in => first_stage_im_out(139),
            re_multiplicator => "0011011011100101", --- 0.857727050781 + j-0.514099121094
            im_multiplicator => "1101111100011001",
            data_re_out => mul_re_out(139),
            data_im_out => mul_im_out(139)
        );

 
    UMUL_140 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(140),
            data_im_in => first_stage_im_out(140),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(140),
            data_im_out => mul_im_out(140)
        );

 
    UMUL_141 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(141),
            data_im_in => first_stage_im_out(141),
            re_multiplicator => "0011001101101000", --- 0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(141),
            data_im_out => mul_im_out(141)
        );

 
    UMUL_142 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(142),
            data_im_in => first_stage_im_out(142),
            re_multiplicator => "0011000101111001", --- 0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(142),
            data_im_out => mul_im_out(142)
        );

 
    UMUL_143 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(143),
            data_im_in => first_stage_im_out(143),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(143),
            data_im_out => mul_im_out(143)
        );

 
    UMUL_144 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(144),
            data_im_in => first_stage_im_out(144),
            re_multiplicator => "0010110101000001", --- 0.707092285156 + j-0.707092285156
            im_multiplicator => "1101001010111111",
            data_re_out => mul_re_out(144),
            data_im_out => mul_im_out(144)
        );

 
    UMUL_145 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(145),
            data_im_in => first_stage_im_out(145),
            re_multiplicator => "0010101011111011", --- 0.671569824219 + j-0.740966796875
            im_multiplicator => "1101000010010100",
            data_re_out => mul_re_out(145),
            data_im_out => mul_im_out(145)
        );

 
    UMUL_146 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(146),
            data_im_in => first_stage_im_out(146),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(146),
            data_im_out => mul_im_out(146)
        );

 
    UMUL_147 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(147),
            data_im_in => first_stage_im_out(147),
            re_multiplicator => "0010011000100000", --- 0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(147),
            data_im_out => mul_im_out(147)
        );

 
    UMUL_148 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(148),
            data_im_in => first_stage_im_out(148),
            re_multiplicator => "0010001110001110", --- 0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(148),
            data_im_out => mul_im_out(148)
        );

 
    UMUL_149 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(149),
            data_im_in => first_stage_im_out(149),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(149),
            data_im_out => mul_im_out(149)
        );

 
    UMUL_150 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(150),
            data_im_in => first_stage_im_out(150),
            re_multiplicator => "0001111000101011", --- 0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(150),
            data_im_out => mul_im_out(150)
        );

 
    UMUL_151 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(151),
            data_im_in => first_stage_im_out(151),
            re_multiplicator => "0001101101011101", --- 0.427551269531 + j-0.903991699219
            im_multiplicator => "1100011000100101",
            data_re_out => mul_re_out(151),
            data_im_out => mul_im_out(151)
        );

 
    UMUL_152 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(152),
            data_im_in => first_stage_im_out(152),
            re_multiplicator => "0001100001111110", --- 0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(152),
            data_im_out => mul_im_out(152)
        );

 
    UMUL_153 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(153),
            data_im_in => first_stage_im_out(153),
            re_multiplicator => "0001010110010000", --- 0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(153),
            data_im_out => mul_im_out(153)
        );

 
    UMUL_154 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(154),
            data_im_in => first_stage_im_out(154),
            re_multiplicator => "0001001010010100", --- 0.290283203125 + j-0.956970214844
            im_multiplicator => "1100001011000001",
            data_re_out => mul_re_out(154),
            data_im_out => mul_im_out(154)
        );

 
    UMUL_155 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(155),
            data_im_in => first_stage_im_out(155),
            re_multiplicator => "0000111110001101", --- 0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(155),
            data_im_out => mul_im_out(155)
        );

 
    UMUL_156 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(156),
            data_im_in => first_stage_im_out(156),
            re_multiplicator => "0000110001111100", --- 0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(156),
            data_im_out => mul_im_out(156)
        );

 
    UMUL_157 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(157),
            data_im_in => first_stage_im_out(157),
            re_multiplicator => "0000100101100100", --- 0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(157),
            data_im_out => mul_im_out(157)
        );

 
    UMUL_158 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(158),
            data_im_in => first_stage_im_out(158),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(158),
            data_im_out => mul_im_out(158)
        );

 
    UMUL_159 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(159),
            data_im_in => first_stage_im_out(159),
            re_multiplicator => "0000001100100100", --- 0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(159),
            data_im_out => mul_im_out(159)
        );

 
    UMUL_160 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(160),
            data_im_in => first_stage_im_out(160),
            data_re_out => mul_re_out(160),
            data_im_out => mul_im_out(160)
        );

 
    UMUL_161 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(161),
            data_im_in => first_stage_im_out(161),
            re_multiplicator => "0011111111100001", --- 0.998107910156 + j-0.0613403320312
            im_multiplicator => "1111110000010011",
            data_re_out => mul_re_out(161),
            data_im_out => mul_im_out(161)
        );

 
    UMUL_162 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(162),
            data_im_in => first_stage_im_out(162),
            re_multiplicator => "0011111110000101", --- 0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(162),
            data_im_out => mul_im_out(162)
        );

 
    UMUL_163 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(163),
            data_im_in => first_stage_im_out(163),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(163),
            data_im_out => mul_im_out(163)
        );

 
    UMUL_164 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(164),
            data_im_in => first_stage_im_out(164),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(164),
            data_im_out => mul_im_out(164)
        );

 
    UMUL_165 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(165),
            data_im_in => first_stage_im_out(165),
            re_multiplicator => "0011110100000011", --- 0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(165),
            data_im_out => mul_im_out(165)
        );

 
    UMUL_166 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(166),
            data_im_in => first_stage_im_out(166),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(166),
            data_im_out => mul_im_out(166)
        );

 
    UMUL_167 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(167),
            data_im_in => first_stage_im_out(167),
            re_multiplicator => "0011101000110000", --- 0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(167),
            data_im_out => mul_im_out(167)
        );

 
    UMUL_168 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(168),
            data_im_in => first_stage_im_out(168),
            re_multiplicator => "0011100001110001", --- 0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(168),
            data_im_out => mul_im_out(168)
        );

 
    UMUL_169 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(169),
            data_im_in => first_stage_im_out(169),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(169),
            data_im_out => mul_im_out(169)
        );

 
    UMUL_170 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(170),
            data_im_in => first_stage_im_out(170),
            re_multiplicator => "0011010001010011", --- 0.817565917969 + j-0.575805664062
            im_multiplicator => "1101101100100110",
            data_re_out => mul_re_out(170),
            data_im_out => mul_im_out(170)
        );

 
    UMUL_171 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(171),
            data_im_in => first_stage_im_out(171),
            re_multiplicator => "0011000111111000", --- 0.78076171875 + j-0.624877929688
            im_multiplicator => "1101100000000010",
            data_re_out => mul_re_out(171),
            data_im_out => mul_im_out(171)
        );

 
    UMUL_172 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(172),
            data_im_in => first_stage_im_out(172),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(172),
            data_im_out => mul_im_out(172)
        );

 
    UMUL_173 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(173),
            data_im_in => first_stage_im_out(173),
            re_multiplicator => "0010110010110010", --- 0.698364257812 + j-0.715759277344
            im_multiplicator => "1101001000110001",
            data_re_out => mul_re_out(173),
            data_im_out => mul_im_out(173)
        );

 
    UMUL_174 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(174),
            data_im_in => first_stage_im_out(174),
            re_multiplicator => "0010100111001110", --- 0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(174),
            data_im_out => mul_im_out(174)
        );

 
    UMUL_175 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(175),
            data_im_in => first_stage_im_out(175),
            re_multiplicator => "0010011011000001", --- 0.605529785156 + j-0.795837402344
            im_multiplicator => "1100110100010001",
            data_re_out => mul_re_out(175),
            data_im_out => mul_im_out(175)
        );

 
    UMUL_176 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(176),
            data_im_in => first_stage_im_out(176),
            re_multiplicator => "0010001110001110", --- 0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(176),
            data_im_out => mul_im_out(176)
        );

 
    UMUL_177 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(177),
            data_im_in => first_stage_im_out(177),
            re_multiplicator => "0010000000111010", --- 0.503540039062 + j-0.863952636719
            im_multiplicator => "1100100010110101",
            data_re_out => mul_re_out(177),
            data_im_out => mul_im_out(177)
        );

 
    UMUL_178 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(178),
            data_im_in => first_stage_im_out(178),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(178),
            data_im_out => mul_im_out(178)
        );

 
    UMUL_179 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(179),
            data_im_in => first_stage_im_out(179),
            re_multiplicator => "0001100100110111", --- 0.393981933594 + j-0.919128417969
            im_multiplicator => "1100010100101101",
            data_re_out => mul_re_out(179),
            data_im_out => mul_im_out(179)
        );

 
    UMUL_180 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(180),
            data_im_in => first_stage_im_out(180),
            re_multiplicator => "0001010110010000", --- 0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(180),
            data_im_out => mul_im_out(180)
        );

 
    UMUL_181 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(181),
            data_im_in => first_stage_im_out(181),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(181),
            data_im_out => mul_im_out(181)
        );

 
    UMUL_182 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(182),
            data_im_in => first_stage_im_out(182),
            re_multiplicator => "0000111000000110", --- 0.219116210938 + j-0.975708007812
            im_multiplicator => "1100000110001110",
            data_re_out => mul_re_out(182),
            data_im_out => mul_im_out(182)
        );

 
    UMUL_183 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(183),
            data_im_in => first_stage_im_out(183),
            re_multiplicator => "0000101000101011", --- 0.158874511719 + j-0.9873046875
            im_multiplicator => "1100000011010000",
            data_re_out => mul_re_out(183),
            data_im_out => mul_im_out(183)
        );

 
    UMUL_184 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(184),
            data_im_in => first_stage_im_out(184),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(184),
            data_im_out => mul_im_out(184)
        );

 
    UMUL_185 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(185),
            data_im_in => first_stage_im_out(185),
            re_multiplicator => "0000001001011011", --- 0.0368041992188 + j-0.999328613281
            im_multiplicator => "1100000000001011",
            data_re_out => mul_re_out(185),
            data_im_out => mul_im_out(185)
        );

 
    UMUL_186 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(186),
            data_im_in => first_stage_im_out(186),
            re_multiplicator => "1111111001101110", --- -0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(186),
            data_im_out => mul_im_out(186)
        );

 
    UMUL_187 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(187),
            data_im_in => first_stage_im_out(187),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(187),
            data_im_out => mul_im_out(187)
        );

 
    UMUL_188 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(188),
            data_im_in => first_stage_im_out(188),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(188),
            data_im_out => mul_im_out(188)
        );

 
    UMUL_189 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(189),
            data_im_in => first_stage_im_out(189),
            re_multiplicator => "1111001010111111", --- -0.207092285156 + j-0.978332519531
            im_multiplicator => "1100000101100011",
            data_re_out => mul_re_out(189),
            data_im_out => mul_im_out(189)
        );

 
    UMUL_190 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(190),
            data_im_in => first_stage_im_out(190),
            re_multiplicator => "1110111011101110", --- -0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(190),
            data_im_out => mul_im_out(190)
        );

 
    UMUL_191 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(191),
            data_im_in => first_stage_im_out(191),
            re_multiplicator => "1110101100101110", --- -0.325317382812 + j-0.945617675781
            im_multiplicator => "1100001101111011",
            data_re_out => mul_re_out(191),
            data_im_out => mul_im_out(191)
        );

 
    UMUL_192 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(192),
            data_im_in => first_stage_im_out(192),
            data_re_out => mul_re_out(192),
            data_im_out => mul_im_out(192)
        );

 
    UMUL_193 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(193),
            data_im_in => first_stage_im_out(193),
            re_multiplicator => "0011111111010100", --- 0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(193),
            data_im_out => mul_im_out(193)
        );

 
    UMUL_194 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(194),
            data_im_in => first_stage_im_out(194),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(194),
            data_im_out => mul_im_out(194)
        );

 
    UMUL_195 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(195),
            data_im_in => first_stage_im_out(195),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(195),
            data_im_out => mul_im_out(195)
        );

 
    UMUL_196 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(196),
            data_im_in => first_stage_im_out(196),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(196),
            data_im_out => mul_im_out(196)
        );

 
    UMUL_197 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(197),
            data_im_in => first_stage_im_out(197),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(197),
            data_im_out => mul_im_out(197)
        );

 
    UMUL_198 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(198),
            data_im_in => first_stage_im_out(198),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(198),
            data_im_out => mul_im_out(198)
        );

 
    UMUL_199 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(199),
            data_im_in => first_stage_im_out(199),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(199),
            data_im_out => mul_im_out(199)
        );

 
    UMUL_200 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(200),
            data_im_in => first_stage_im_out(200),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(200),
            data_im_out => mul_im_out(200)
        );

 
    UMUL_201 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(201),
            data_im_in => first_stage_im_out(201),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(201),
            data_im_out => mul_im_out(201)
        );

 
    UMUL_202 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(202),
            data_im_in => first_stage_im_out(202),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(202),
            data_im_out => mul_im_out(202)
        );

 
    UMUL_203 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(203),
            data_im_in => first_stage_im_out(203),
            re_multiplicator => "0010110000100001", --- 0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(203),
            data_im_out => mul_im_out(203)
        );

 
    UMUL_204 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(204),
            data_im_in => first_stage_im_out(204),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(204),
            data_im_out => mul_im_out(204)
        );

 
    UMUL_205 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(205),
            data_im_in => first_stage_im_out(205),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j-0.817565917969
            im_multiplicator => "1100101110101101",
            data_re_out => mul_re_out(205),
            data_im_out => mul_im_out(205)
        );

 
    UMUL_206 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(206),
            data_im_in => first_stage_im_out(206),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(206),
            data_im_out => mul_im_out(206)
        );

 
    UMUL_207 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(207),
            data_im_in => first_stage_im_out(207),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(207),
            data_im_out => mul_im_out(207)
        );

 
    UMUL_208 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(208),
            data_im_in => first_stage_im_out(208),
            re_multiplicator => "0001100001111110", --- 0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(208),
            data_im_out => mul_im_out(208)
        );

 
    UMUL_209 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(209),
            data_im_in => first_stage_im_out(209),
            re_multiplicator => "0001010000010011", --- 0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(209),
            data_im_out => mul_im_out(209)
        );

 
    UMUL_210 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(210),
            data_im_in => first_stage_im_out(210),
            re_multiplicator => "0000111110001101", --- 0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(210),
            data_im_out => mul_im_out(210)
        );

 
    UMUL_211 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(211),
            data_im_in => first_stage_im_out(211),
            re_multiplicator => "0000101011110001", --- 0.170959472656 + j-0.985290527344
            im_multiplicator => "1100000011110001",
            data_re_out => mul_re_out(211),
            data_im_out => mul_im_out(211)
        );

 
    UMUL_212 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(212),
            data_im_in => first_stage_im_out(212),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(212),
            data_im_out => mul_im_out(212)
        );

 
    UMUL_213 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(213),
            data_im_in => first_stage_im_out(213),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(213),
            data_im_out => mul_im_out(213)
        );

 
    UMUL_214 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(214),
            data_im_in => first_stage_im_out(214),
            re_multiplicator => "1111110011011100", --- -0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(214),
            data_im_out => mul_im_out(214)
        );

 
    UMUL_215 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(215),
            data_im_in => first_stage_im_out(215),
            re_multiplicator => "1111100000101010", --- -0.122436523438 + j-0.992492675781
            im_multiplicator => "1100000001111011",
            data_re_out => mul_re_out(215),
            data_im_out => mul_im_out(215)
        );

 
    UMUL_216 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(216),
            data_im_in => first_stage_im_out(216),
            re_multiplicator => "1111001110000100", --- -0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(216),
            data_im_out => mul_im_out(216)
        );

 
    UMUL_217 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(217),
            data_im_in => first_stage_im_out(217),
            re_multiplicator => "1110111011101110", --- -0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(217),
            data_im_out => mul_im_out(217)
        );

 
    UMUL_218 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(218),
            data_im_in => first_stage_im_out(218),
            re_multiplicator => "1110101001110000", --- -0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(218),
            data_im_out => mul_im_out(218)
        );

 
    UMUL_219 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(219),
            data_im_in => first_stage_im_out(219),
            re_multiplicator => "1110011000010001", --- -0.405212402344 + j-0.914184570312
            im_multiplicator => "1100010101111110",
            data_re_out => mul_re_out(219),
            data_im_out => mul_im_out(219)
        );

 
    UMUL_220 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(220),
            data_im_in => first_stage_im_out(220),
            re_multiplicator => "1110000111010101", --- -0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(220),
            data_im_out => mul_im_out(220)
        );

 
    UMUL_221 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(221),
            data_im_in => first_stage_im_out(221),
            re_multiplicator => "1101110111000011", --- -0.534973144531 + j-0.844848632812
            im_multiplicator => "1100100111101110",
            data_re_out => mul_re_out(221),
            data_im_out => mul_im_out(221)
        );

 
    UMUL_222 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(222),
            data_im_in => first_stage_im_out(222),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(222),
            data_im_out => mul_im_out(222)
        );

 
    UMUL_223 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(223),
            data_im_in => first_stage_im_out(223),
            re_multiplicator => "1101011000110010", --- -0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(223),
            data_im_out => mul_im_out(223)
        );

 
    UMUL_224 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(224),
            data_im_in => first_stage_im_out(224),
            data_re_out => mul_re_out(224),
            data_im_out => mul_im_out(224)
        );

 
    UMUL_225 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(225),
            data_im_in => first_stage_im_out(225),
            re_multiplicator => "0011111111000100", --- 0.996337890625 + j-0.0858154296875
            im_multiplicator => "1111101010000010",
            data_re_out => mul_re_out(225),
            data_im_out => mul_im_out(225)
        );

 
    UMUL_226 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(226),
            data_im_in => first_stage_im_out(226),
            re_multiplicator => "0011111100001111", --- 0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(226),
            data_im_out => mul_im_out(226)
        );

 
    UMUL_227 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(227),
            data_im_in => first_stage_im_out(227),
            re_multiplicator => "0011110111100011", --- 0.966979980469 + j-0.2548828125
            im_multiplicator => "1110111110110000",
            data_re_out => mul_re_out(227),
            data_im_out => mul_im_out(227)
        );

 
    UMUL_228 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(228),
            data_im_in => first_stage_im_out(228),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(228),
            data_im_out => mul_im_out(228)
        );

 
    UMUL_229 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(229),
            data_im_in => first_stage_im_out(229),
            re_multiplicator => "0011101000110000", --- 0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(229),
            data_im_out => mul_im_out(229)
        );

 
    UMUL_230 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(230),
            data_im_in => first_stage_im_out(230),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(230),
            data_im_out => mul_im_out(230)
        );

 
    UMUL_231 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(231),
            data_im_in => first_stage_im_out(231),
            re_multiplicator => "0011010011000110", --- 0.824584960938 + j-0.565734863281
            im_multiplicator => "1101101111001011",
            data_re_out => mul_re_out(231),
            data_im_out => mul_im_out(231)
        );

 
    UMUL_232 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(232),
            data_im_in => first_stage_im_out(232),
            re_multiplicator => "0011000101111001", --- 0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(232),
            data_im_out => mul_im_out(232)
        );

 
    UMUL_233 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(233),
            data_im_in => first_stage_im_out(233),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(233),
            data_im_out => mul_im_out(233)
        );

 
    UMUL_234 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(234),
            data_im_in => first_stage_im_out(234),
            re_multiplicator => "0010100111001110", --- 0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(234),
            data_im_out => mul_im_out(234)
        );

 
    UMUL_235 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(235),
            data_im_in => first_stage_im_out(235),
            re_multiplicator => "0010010101111110", --- 0.585815429688 + j-0.810485839844
            im_multiplicator => "1100110000100001",
            data_re_out => mul_re_out(235),
            data_im_out => mul_im_out(235)
        );

 
    UMUL_236 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(236),
            data_im_in => first_stage_im_out(236),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(236),
            data_im_out => mul_im_out(236)
        );

 
    UMUL_237 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(237),
            data_im_in => first_stage_im_out(237),
            re_multiplicator => "0001110000010010", --- 0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(237),
            data_im_out => mul_im_out(237)
        );

 
    UMUL_238 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(238),
            data_im_in => first_stage_im_out(238),
            re_multiplicator => "0001011100001001", --- 0.359924316406 + j-0.932983398438
            im_multiplicator => "1100010001001010",
            data_re_out => mul_re_out(238),
            data_im_out => mul_im_out(238)
        );

 
    UMUL_239 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(239),
            data_im_in => first_stage_im_out(239),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(239),
            data_im_out => mul_im_out(239)
        );

 
    UMUL_240 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(240),
            data_im_in => first_stage_im_out(240),
            re_multiplicator => "0000110001111100", --- 0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(240),
            data_im_out => mul_im_out(240)
        );

 
    UMUL_241 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(241),
            data_im_in => first_stage_im_out(241),
            re_multiplicator => "0000011100001110", --- 0.110229492188 + j-0.993896484375
            im_multiplicator => "1100000001100100",
            data_re_out => mul_re_out(241),
            data_im_out => mul_im_out(241)
        );

 
    UMUL_242 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(242),
            data_im_in => first_stage_im_out(242),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(242),
            data_im_out => mul_im_out(242)
        );

 
    UMUL_243 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(243),
            data_im_in => first_stage_im_out(243),
            re_multiplicator => "1111110000010011", --- -0.0613403320312 + j-0.998107910156
            im_multiplicator => "1100000000011111",
            data_re_out => mul_re_out(243),
            data_im_out => mul_im_out(243)
        );

 
    UMUL_244 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(244),
            data_im_in => first_stage_im_out(244),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(244),
            data_im_out => mul_im_out(244)
        );

 
    UMUL_245 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(245),
            data_im_in => first_stage_im_out(245),
            re_multiplicator => "1111000100110110", --- -0.231079101562 + j-0.972961425781
            im_multiplicator => "1100000110111011",
            data_re_out => mul_re_out(245),
            data_im_out => mul_im_out(245)
        );

 
    UMUL_246 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(246),
            data_im_in => first_stage_im_out(246),
            re_multiplicator => "1110101111101101", --- -0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(246),
            data_im_out => mul_im_out(246)
        );

 
    UMUL_247 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(247),
            data_im_in => first_stage_im_out(247),
            re_multiplicator => "1110011011001001", --- -0.393981933594 + j-0.919128417969
            im_multiplicator => "1100010100101101",
            data_re_out => mul_re_out(247),
            data_im_out => mul_im_out(247)
        );

 
    UMUL_248 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(248),
            data_im_in => first_stage_im_out(248),
            re_multiplicator => "1110000111010101", --- -0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(248),
            data_im_out => mul_im_out(248)
        );

 
    UMUL_249 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(249),
            data_im_in => first_stage_im_out(249),
            re_multiplicator => "1101110100011001", --- -0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(249),
            data_im_out => mul_im_out(249)
        );

 
    UMUL_250 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(250),
            data_im_in => first_stage_im_out(250),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j-0.788330078125
            im_multiplicator => "1100110110001100",
            data_re_out => mul_re_out(250),
            data_im_out => mul_im_out(250)
        );

 
    UMUL_251 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(251),
            data_im_in => first_stage_im_out(251),
            re_multiplicator => "1101010001110001", --- -0.680603027344 + j-0.732666015625
            im_multiplicator => "1101000100011100",
            data_re_out => mul_re_out(251),
            data_im_out => mul_im_out(251)
        );

 
    UMUL_252 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(252),
            data_im_in => first_stage_im_out(252),
            re_multiplicator => "1101000010010100", --- -0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(252),
            data_im_out => mul_im_out(252)
        );

 
    UMUL_253 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(253),
            data_im_in => first_stage_im_out(253),
            re_multiplicator => "1100110100010001", --- -0.795837402344 + j-0.605529785156
            im_multiplicator => "1101100100111111",
            data_re_out => mul_re_out(253),
            data_im_out => mul_im_out(253)
        );

 
    UMUL_254 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(254),
            data_im_in => first_stage_im_out(254),
            re_multiplicator => "1100100111101110", --- -0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(254),
            data_im_out => mul_im_out(254)
        );

 
    UMUL_255 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(255),
            data_im_in => first_stage_im_out(255),
            re_multiplicator => "1100011100110001", --- -0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(255),
            data_im_out => mul_im_out(255)
        );

 
    UMUL_256 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(256),
            data_im_in => first_stage_im_out(256),
            data_re_out => mul_re_out(256),
            data_im_out => mul_im_out(256)
        );

 
    UMUL_257 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(257),
            data_im_in => first_stage_im_out(257),
            re_multiplicator => "0011111110110001", --- 0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(257),
            data_im_out => mul_im_out(257)
        );

 
    UMUL_258 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(258),
            data_im_in => first_stage_im_out(258),
            re_multiplicator => "0011111011000101", --- 0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(258),
            data_im_out => mul_im_out(258)
        );

 
    UMUL_259 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(259),
            data_im_in => first_stage_im_out(259),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(259),
            data_im_out => mul_im_out(259)
        );

 
    UMUL_260 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(260),
            data_im_in => first_stage_im_out(260),
            re_multiplicator => "0011101100100001", --- 0.923889160156 + j-0.382690429688
            im_multiplicator => "1110011110000010",
            data_re_out => mul_re_out(260),
            data_im_out => mul_im_out(260)
        );

 
    UMUL_261 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(261),
            data_im_in => first_stage_im_out(261),
            re_multiplicator => "0011100001110001", --- 0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(261),
            data_im_out => mul_im_out(261)
        );

 
    UMUL_262 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(262),
            data_im_in => first_stage_im_out(262),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(262),
            data_im_out => mul_im_out(262)
        );

 
    UMUL_263 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(263),
            data_im_in => first_stage_im_out(263),
            re_multiplicator => "0011000101111001", --- 0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(263),
            data_im_out => mul_im_out(263)
        );

 
    UMUL_264 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(264),
            data_im_in => first_stage_im_out(264),
            re_multiplicator => "0010110101000001", --- 0.707092285156 + j-0.707092285156
            im_multiplicator => "1101001010111111",
            data_re_out => mul_re_out(264),
            data_im_out => mul_im_out(264)
        );

 
    UMUL_265 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(265),
            data_im_in => first_stage_im_out(265),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(265),
            data_im_out => mul_im_out(265)
        );

 
    UMUL_266 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(266),
            data_im_in => first_stage_im_out(266),
            re_multiplicator => "0010001110001110", --- 0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(266),
            data_im_out => mul_im_out(266)
        );

 
    UMUL_267 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(267),
            data_im_in => first_stage_im_out(267),
            re_multiplicator => "0001111000101011", --- 0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(267),
            data_im_out => mul_im_out(267)
        );

 
    UMUL_268 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(268),
            data_im_in => first_stage_im_out(268),
            re_multiplicator => "0001100001111110", --- 0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(268),
            data_im_out => mul_im_out(268)
        );

 
    UMUL_269 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(269),
            data_im_in => first_stage_im_out(269),
            re_multiplicator => "0001001010010100", --- 0.290283203125 + j-0.956970214844
            im_multiplicator => "1100001011000001",
            data_re_out => mul_re_out(269),
            data_im_out => mul_im_out(269)
        );

 
    UMUL_270 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(270),
            data_im_in => first_stage_im_out(270),
            re_multiplicator => "0000110001111100", --- 0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(270),
            data_im_out => mul_im_out(270)
        );

 
    UMUL_271 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(271),
            data_im_in => first_stage_im_out(271),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(271),
            data_im_out => mul_im_out(271)
        );

 
    UMUL_272 : multiplier_mulminusj
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(272),
            data_im_in => first_stage_im_out(272),
            data_re_out => mul_re_out(272),
            data_im_out => mul_im_out(272)
        );

 
    UMUL_273 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(273),
            data_im_in => first_stage_im_out(273),
            re_multiplicator => "1111100110111010", --- -0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(273),
            data_im_out => mul_im_out(273)
        );

 
    UMUL_274 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(274),
            data_im_in => first_stage_im_out(274),
            re_multiplicator => "1111001110000100", --- -0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(274),
            data_im_out => mul_im_out(274)
        );

 
    UMUL_275 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(275),
            data_im_in => first_stage_im_out(275),
            re_multiplicator => "1110110101101100", --- -0.290283203125 + j-0.956970214844
            im_multiplicator => "1100001011000001",
            data_re_out => mul_re_out(275),
            data_im_out => mul_im_out(275)
        );

 
    UMUL_276 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(276),
            data_im_in => first_stage_im_out(276),
            re_multiplicator => "1110011110000010", --- -0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(276),
            data_im_out => mul_im_out(276)
        );

 
    UMUL_277 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(277),
            data_im_in => first_stage_im_out(277),
            re_multiplicator => "1110000111010101", --- -0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(277),
            data_im_out => mul_im_out(277)
        );

 
    UMUL_278 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(278),
            data_im_in => first_stage_im_out(278),
            re_multiplicator => "1101110001110010", --- -0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(278),
            data_im_out => mul_im_out(278)
        );

 
    UMUL_279 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(279),
            data_im_in => first_stage_im_out(279),
            re_multiplicator => "1101011101100110", --- -0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(279),
            data_im_out => mul_im_out(279)
        );

 
    UMUL_280 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(280),
            data_im_in => first_stage_im_out(280),
            re_multiplicator => "1101001010111111", --- -0.707092285156 + j-0.707092285156
            im_multiplicator => "1101001010111111",
            data_re_out => mul_re_out(280),
            data_im_out => mul_im_out(280)
        );

 
    UMUL_281 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(281),
            data_im_in => first_stage_im_out(281),
            re_multiplicator => "1100111010000111", --- -0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(281),
            data_im_out => mul_im_out(281)
        );

 
    UMUL_282 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(282),
            data_im_in => first_stage_im_out(282),
            re_multiplicator => "1100101011001001", --- -0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(282),
            data_im_out => mul_im_out(282)
        );

 
    UMUL_283 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(283),
            data_im_in => first_stage_im_out(283),
            re_multiplicator => "1100011110001111", --- -0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(283),
            data_im_out => mul_im_out(283)
        );

 
    UMUL_284 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(284),
            data_im_in => first_stage_im_out(284),
            re_multiplicator => "1100010011011111", --- -0.923889160156 + j-0.382690429688
            im_multiplicator => "1110011110000010",
            data_re_out => mul_re_out(284),
            data_im_out => mul_im_out(284)
        );

 
    UMUL_285 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(285),
            data_im_in => first_stage_im_out(285),
            re_multiplicator => "1100001011000001", --- -0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(285),
            data_im_out => mul_im_out(285)
        );

 
    UMUL_286 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(286),
            data_im_in => first_stage_im_out(286),
            re_multiplicator => "1100000100111011", --- -0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(286),
            data_im_out => mul_im_out(286)
        );

 
    UMUL_287 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(287),
            data_im_in => first_stage_im_out(287),
            re_multiplicator => "1100000001001111", --- -0.995178222656 + j-0.0980224609375
            im_multiplicator => "1111100110111010",
            data_re_out => mul_re_out(287),
            data_im_out => mul_im_out(287)
        );

 
    UMUL_288 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(288),
            data_im_in => first_stage_im_out(288),
            data_re_out => mul_re_out(288),
            data_im_out => mul_im_out(288)
        );

 
    UMUL_289 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(289),
            data_im_in => first_stage_im_out(289),
            re_multiplicator => "0011111110011100", --- 0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(289),
            data_im_out => mul_im_out(289)
        );

 
    UMUL_290 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(290),
            data_im_in => first_stage_im_out(290),
            re_multiplicator => "0011111001110010", --- 0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(290),
            data_im_out => mul_im_out(290)
        );

 
    UMUL_291 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(291),
            data_im_in => first_stage_im_out(291),
            re_multiplicator => "0011110010000101", --- 0.945617675781 + j-0.325317382812
            im_multiplicator => "1110101100101110",
            data_re_out => mul_re_out(291),
            data_im_out => mul_im_out(291)
        );

 
    UMUL_292 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(292),
            data_im_in => first_stage_im_out(292),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(292),
            data_im_out => mul_im_out(292)
        );

 
    UMUL_293 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(293),
            data_im_in => first_stage_im_out(293),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(293),
            data_im_out => mul_im_out(293)
        );

 
    UMUL_294 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(294),
            data_im_in => first_stage_im_out(294),
            re_multiplicator => "0011001001110100", --- 0.788330078125 + j-0.615234375
            im_multiplicator => "1101100010100000",
            data_re_out => mul_re_out(294),
            data_im_out => mul_im_out(294)
        );

 
    UMUL_295 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(295),
            data_im_in => first_stage_im_out(295),
            re_multiplicator => "0010110111001111", --- 0.715759277344 + j-0.698364257812
            im_multiplicator => "1101001101001110",
            data_re_out => mul_re_out(295),
            data_im_out => mul_im_out(295)
        );

 
    UMUL_296 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(296),
            data_im_in => first_stage_im_out(296),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(296),
            data_im_out => mul_im_out(296)
        );

 
    UMUL_297 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(297),
            data_im_in => first_stage_im_out(297),
            re_multiplicator => "0010001011100111", --- 0.545349121094 + j-0.838195800781
            im_multiplicator => "1100101001011011",
            data_re_out => mul_re_out(297),
            data_im_out => mul_im_out(297)
        );

 
    UMUL_298 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(298),
            data_im_in => first_stage_im_out(298),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(298),
            data_im_out => mul_im_out(298)
        );

 
    UMUL_299 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(299),
            data_im_in => first_stage_im_out(299),
            re_multiplicator => "0001011001001100", --- 0.348388671875 + j-0.937316894531
            im_multiplicator => "1100010000000011",
            data_re_out => mul_re_out(299),
            data_im_out => mul_im_out(299)
        );

 
    UMUL_300 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(300),
            data_im_in => first_stage_im_out(300),
            re_multiplicator => "0000111110001101", --- 0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(300),
            data_im_out => mul_im_out(300)
        );

 
    UMUL_301 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(301),
            data_im_in => first_stage_im_out(301),
            re_multiplicator => "0000100010011101", --- 0.134582519531 + j-0.990905761719
            im_multiplicator => "1100000010010101",
            data_re_out => mul_re_out(301),
            data_im_out => mul_im_out(301)
        );

 
    UMUL_302 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(302),
            data_im_in => first_stage_im_out(302),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(302),
            data_im_out => mul_im_out(302)
        );

 
    UMUL_303 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(303),
            data_im_in => first_stage_im_out(303),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(303),
            data_im_out => mul_im_out(303)
        );

 
    UMUL_304 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(304),
            data_im_in => first_stage_im_out(304),
            re_multiplicator => "1111001110000100", --- -0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(304),
            data_im_out => mul_im_out(304)
        );

 
    UMUL_305 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(305),
            data_im_in => first_stage_im_out(305),
            re_multiplicator => "1110110010101100", --- -0.302001953125 + j-0.953308105469
            im_multiplicator => "1100001011111101",
            data_re_out => mul_re_out(305),
            data_im_out => mul_im_out(305)
        );

 
    UMUL_306 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(306),
            data_im_in => first_stage_im_out(306),
            re_multiplicator => "1110011000010001", --- -0.405212402344 + j-0.914184570312
            im_multiplicator => "1100010101111110",
            data_re_out => mul_re_out(306),
            data_im_out => mul_im_out(306)
        );

 
    UMUL_307 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(307),
            data_im_in => first_stage_im_out(307),
            re_multiplicator => "1101111111000110", --- -0.503540039062 + j-0.863952636719
            im_multiplicator => "1100100010110101",
            data_re_out => mul_re_out(307),
            data_im_out => mul_im_out(307)
        );

 
    UMUL_308 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(308),
            data_im_in => first_stage_im_out(308),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(308),
            data_im_out => mul_im_out(308)
        );

 
    UMUL_309 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(309),
            data_im_in => first_stage_im_out(309),
            re_multiplicator => "1101010001110001", --- -0.680603027344 + j-0.732666015625
            im_multiplicator => "1101000100011100",
            data_re_out => mul_re_out(309),
            data_im_out => mul_im_out(309)
        );

 
    UMUL_310 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(310),
            data_im_in => first_stage_im_out(310),
            re_multiplicator => "1100111110001010", --- -0.757202148438 + j-0.653198242188
            im_multiplicator => "1101011000110010",
            data_re_out => mul_re_out(310),
            data_im_out => mul_im_out(310)
        );

 
    UMUL_311 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(311),
            data_im_in => first_stage_im_out(311),
            re_multiplicator => "1100101100111010", --- -0.824584960938 + j-0.565734863281
            im_multiplicator => "1101101111001011",
            data_re_out => mul_re_out(311),
            data_im_out => mul_im_out(311)
        );

 
    UMUL_312 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(312),
            data_im_in => first_stage_im_out(312),
            re_multiplicator => "1100011110001111", --- -0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(312),
            data_im_out => mul_im_out(312)
        );

 
    UMUL_313 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(313),
            data_im_in => first_stage_im_out(313),
            re_multiplicator => "1100010010010011", --- -0.928527832031 + j-0.371337890625
            im_multiplicator => "1110100000111100",
            data_re_out => mul_re_out(313),
            data_im_out => mul_im_out(313)
        );

 
    UMUL_314 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(314),
            data_im_in => first_stage_im_out(314),
            re_multiplicator => "1100001001010001", --- -0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(314),
            data_im_out => mul_im_out(314)
        );

 
    UMUL_315 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(315),
            data_im_in => first_stage_im_out(315),
            re_multiplicator => "1100000011010000", --- -0.9873046875 + j-0.158874511719
            im_multiplicator => "1111010111010101",
            data_re_out => mul_re_out(315),
            data_im_out => mul_im_out(315)
        );

 
    UMUL_316 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(316),
            data_im_in => first_stage_im_out(316),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(316),
            data_im_out => mul_im_out(316)
        );

 
    UMUL_317 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(317),
            data_im_in => first_stage_im_out(317),
            re_multiplicator => "1100000000011111", --- -0.998107910156 + j0.0613403320312
            im_multiplicator => "0000001111101101",
            data_re_out => mul_re_out(317),
            data_im_out => mul_im_out(317)
        );

 
    UMUL_318 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(318),
            data_im_in => first_stage_im_out(318),
            re_multiplicator => "1100000011110001", --- -0.985290527344 + j0.170959472656
            im_multiplicator => "0000101011110001",
            data_re_out => mul_re_out(318),
            data_im_out => mul_im_out(318)
        );

 
    UMUL_319 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(319),
            data_im_in => first_stage_im_out(319),
            re_multiplicator => "1100001010001000", --- -0.96044921875 + j0.278503417969
            im_multiplicator => "0001000111010011",
            data_re_out => mul_re_out(319),
            data_im_out => mul_im_out(319)
        );

 
    UMUL_320 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(320),
            data_im_in => first_stage_im_out(320),
            data_re_out => mul_re_out(320),
            data_im_out => mul_im_out(320)
        );

 
    UMUL_321 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(321),
            data_im_in => first_stage_im_out(321),
            re_multiplicator => "0011111110000101", --- 0.992492675781 + j-0.122436523438
            im_multiplicator => "1111100000101010",
            data_re_out => mul_re_out(321),
            data_im_out => mul_im_out(321)
        );

 
    UMUL_322 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(322),
            data_im_in => first_stage_im_out(322),
            re_multiplicator => "0011111000010101", --- 0.970031738281 + j-0.242980957031
            im_multiplicator => "1111000001110011",
            data_re_out => mul_re_out(322),
            data_im_out => mul_im_out(322)
        );

 
    UMUL_323 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(323),
            data_im_in => first_stage_im_out(323),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(323),
            data_im_out => mul_im_out(323)
        );

 
    UMUL_324 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(324),
            data_im_in => first_stage_im_out(324),
            re_multiplicator => "0011100001110001", --- 0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(324),
            data_im_out => mul_im_out(324)
        );

 
    UMUL_325 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(325),
            data_im_in => first_stage_im_out(325),
            re_multiplicator => "0011010001010011", --- 0.817565917969 + j-0.575805664062
            im_multiplicator => "1101101100100110",
            data_re_out => mul_re_out(325),
            data_im_out => mul_im_out(325)
        );

 
    UMUL_326 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(326),
            data_im_in => first_stage_im_out(326),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(326),
            data_im_out => mul_im_out(326)
        );

 
    UMUL_327 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(327),
            data_im_in => first_stage_im_out(327),
            re_multiplicator => "0010100111001110", --- 0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(327),
            data_im_out => mul_im_out(327)
        );

 
    UMUL_328 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(328),
            data_im_in => first_stage_im_out(328),
            re_multiplicator => "0010001110001110", --- 0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(328),
            data_im_out => mul_im_out(328)
        );

 
    UMUL_329 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(329),
            data_im_in => first_stage_im_out(329),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(329),
            data_im_out => mul_im_out(329)
        );

 
    UMUL_330 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(330),
            data_im_in => first_stage_im_out(330),
            re_multiplicator => "0001010110010000", --- 0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(330),
            data_im_out => mul_im_out(330)
        );

 
    UMUL_331 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(331),
            data_im_in => first_stage_im_out(331),
            re_multiplicator => "0000111000000110", --- 0.219116210938 + j-0.975708007812
            im_multiplicator => "1100000110001110",
            data_re_out => mul_re_out(331),
            data_im_out => mul_im_out(331)
        );

 
    UMUL_332 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(332),
            data_im_in => first_stage_im_out(332),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(332),
            data_im_out => mul_im_out(332)
        );

 
    UMUL_333 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(333),
            data_im_in => first_stage_im_out(333),
            re_multiplicator => "1111111001101110", --- -0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(333),
            data_im_out => mul_im_out(333)
        );

 
    UMUL_334 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(334),
            data_im_in => first_stage_im_out(334),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(334),
            data_im_out => mul_im_out(334)
        );

 
    UMUL_335 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(335),
            data_im_in => first_stage_im_out(335),
            re_multiplicator => "1110111011101110", --- -0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(335),
            data_im_out => mul_im_out(335)
        );

 
    UMUL_336 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(336),
            data_im_in => first_stage_im_out(336),
            re_multiplicator => "1110011110000010", --- -0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(336),
            data_im_out => mul_im_out(336)
        );

 
    UMUL_337 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(337),
            data_im_in => first_stage_im_out(337),
            re_multiplicator => "1110000001110100", --- -0.492919921875 + j-0.8701171875
            im_multiplicator => "1100100001010000",
            data_re_out => mul_re_out(337),
            data_im_out => mul_im_out(337)
        );

 
    UMUL_338 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(338),
            data_im_in => first_stage_im_out(338),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(338),
            data_im_out => mul_im_out(338)
        );

 
    UMUL_339 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(339),
            data_im_in => first_stage_im_out(339),
            re_multiplicator => "1101001111011111", --- -0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(339),
            data_im_out => mul_im_out(339)
        );

 
    UMUL_340 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(340),
            data_im_in => first_stage_im_out(340),
            re_multiplicator => "1100111010000111", --- -0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(340),
            data_im_out => mul_im_out(340)
        );

 
    UMUL_341 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(341),
            data_im_in => first_stage_im_out(341),
            re_multiplicator => "1100100111101110", --- -0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(341),
            data_im_out => mul_im_out(341)
        );

 
    UMUL_342 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(342),
            data_im_in => first_stage_im_out(342),
            re_multiplicator => "1100011000100101", --- -0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(342),
            data_im_out => mul_im_out(342)
        );

 
    UMUL_343 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(343),
            data_im_in => first_stage_im_out(343),
            re_multiplicator => "1100001100111011", --- -0.949523925781 + j-0.313659667969
            im_multiplicator => "1110101111101101",
            data_re_out => mul_re_out(343),
            data_im_out => mul_im_out(343)
        );

 
    UMUL_344 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(344),
            data_im_in => first_stage_im_out(344),
            re_multiplicator => "1100000100111011", --- -0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(344),
            data_im_out => mul_im_out(344)
        );

 
    UMUL_345 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(345),
            data_im_in => first_stage_im_out(345),
            re_multiplicator => "1100000000101100", --- -0.997314453125 + j-0.0735473632812
            im_multiplicator => "1111101101001011",
            data_re_out => mul_re_out(345),
            data_im_out => mul_im_out(345)
        );

 
    UMUL_346 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(346),
            data_im_in => first_stage_im_out(346),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j0.049072265625
            im_multiplicator => "0000001100100100",
            data_re_out => mul_re_out(346),
            data_im_out => mul_im_out(346)
        );

 
    UMUL_347 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(347),
            data_im_in => first_stage_im_out(347),
            re_multiplicator => "1100000011110001", --- -0.985290527344 + j0.170959472656
            im_multiplicator => "0000101011110001",
            data_re_out => mul_re_out(347),
            data_im_out => mul_im_out(347)
        );

 
    UMUL_348 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(348),
            data_im_in => first_stage_im_out(348),
            re_multiplicator => "1100001011000001", --- -0.956970214844 + j0.290283203125
            im_multiplicator => "0001001010010100",
            data_re_out => mul_re_out(348),
            data_im_out => mul_im_out(348)
        );

 
    UMUL_349 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(349),
            data_im_in => first_stage_im_out(349),
            re_multiplicator => "1100010101111110", --- -0.914184570312 + j0.405212402344
            im_multiplicator => "0001100111101111",
            data_re_out => mul_re_out(349),
            data_im_out => mul_im_out(349)
        );

 
    UMUL_350 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(350),
            data_im_in => first_stage_im_out(350),
            re_multiplicator => "1100100100011011", --- -0.857727050781 + j0.514099121094
            im_multiplicator => "0010000011100111",
            data_re_out => mul_re_out(350),
            data_im_out => mul_im_out(350)
        );

 
    UMUL_351 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(351),
            data_im_in => first_stage_im_out(351),
            re_multiplicator => "1100110110001100", --- -0.788330078125 + j0.615234375
            im_multiplicator => "0010011101100000",
            data_re_out => mul_re_out(351),
            data_im_out => mul_im_out(351)
        );

 
    UMUL_352 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(352),
            data_im_in => first_stage_im_out(352),
            data_re_out => mul_re_out(352),
            data_im_out => mul_im_out(352)
        );

 
    UMUL_353 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(353),
            data_im_in => first_stage_im_out(353),
            re_multiplicator => "0011111101101011", --- 0.990905761719 + j-0.134582519531
            im_multiplicator => "1111011101100011",
            data_re_out => mul_re_out(353),
            data_im_out => mul_im_out(353)
        );

 
    UMUL_354 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(354),
            data_im_in => first_stage_im_out(354),
            re_multiplicator => "0011110110101111", --- 0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(354),
            data_im_out => mul_im_out(354)
        );

 
    UMUL_355 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(355),
            data_im_in => first_stage_im_out(355),
            re_multiplicator => "0011101011010011", --- 0.919128417969 + j-0.393981933594
            im_multiplicator => "1110011011001001",
            data_re_out => mul_re_out(355),
            data_im_out => mul_im_out(355)
        );

 
    UMUL_356 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(356),
            data_im_in => first_stage_im_out(356),
            re_multiplicator => "0011011011100101", --- 0.857727050781 + j-0.514099121094
            im_multiplicator => "1101111100011001",
            data_re_out => mul_re_out(356),
            data_im_out => mul_im_out(356)
        );

 
    UMUL_357 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(357),
            data_im_in => first_stage_im_out(357),
            re_multiplicator => "0011000111111000", --- 0.78076171875 + j-0.624877929688
            im_multiplicator => "1101100000000010",
            data_re_out => mul_re_out(357),
            data_im_out => mul_im_out(357)
        );

 
    UMUL_358 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(358),
            data_im_in => first_stage_im_out(358),
            re_multiplicator => "0010110000100001", --- 0.689514160156 + j-0.724243164062
            im_multiplicator => "1101000110100110",
            data_re_out => mul_re_out(358),
            data_im_out => mul_im_out(358)
        );

 
    UMUL_359 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(359),
            data_im_in => first_stage_im_out(359),
            re_multiplicator => "0010010101111110", --- 0.585815429688 + j-0.810485839844
            im_multiplicator => "1100110000100001",
            data_re_out => mul_re_out(359),
            data_im_out => mul_im_out(359)
        );

 
    UMUL_360 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(360),
            data_im_in => first_stage_im_out(360),
            re_multiplicator => "0001111000101011", --- 0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(360),
            data_im_out => mul_im_out(360)
        );

 
    UMUL_361 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(361),
            data_im_in => first_stage_im_out(361),
            re_multiplicator => "0001011001001100", --- 0.348388671875 + j-0.937316894531
            im_multiplicator => "1100010000000011",
            data_re_out => mul_re_out(361),
            data_im_out => mul_im_out(361)
        );

 
    UMUL_362 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(362),
            data_im_in => first_stage_im_out(362),
            re_multiplicator => "0000111000000110", --- 0.219116210938 + j-0.975708007812
            im_multiplicator => "1100000110001110",
            data_re_out => mul_re_out(362),
            data_im_out => mul_im_out(362)
        );

 
    UMUL_363 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(363),
            data_im_in => first_stage_im_out(363),
            re_multiplicator => "0000010101111110", --- 0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(363),
            data_im_out => mul_im_out(363)
        );

 
    UMUL_364 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(364),
            data_im_in => first_stage_im_out(364),
            re_multiplicator => "1111110011011100", --- -0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(364),
            data_im_out => mul_im_out(364)
        );

 
    UMUL_365 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(365),
            data_im_in => first_stage_im_out(365),
            re_multiplicator => "1111010001001001", --- -0.183044433594 + j-0.983093261719
            im_multiplicator => "1100000100010101",
            data_re_out => mul_re_out(365),
            data_im_out => mul_im_out(365)
        );

 
    UMUL_366 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(366),
            data_im_in => first_stage_im_out(366),
            re_multiplicator => "1110101111101101", --- -0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(366),
            data_im_out => mul_im_out(366)
        );

 
    UMUL_367 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(367),
            data_im_in => first_stage_im_out(367),
            re_multiplicator => "1110001111101110", --- -0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(367),
            data_im_out => mul_im_out(367)
        );

 
    UMUL_368 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(368),
            data_im_in => first_stage_im_out(368),
            re_multiplicator => "1101110001110010", --- -0.555541992188 + j-0.831481933594
            im_multiplicator => "1100101011001001",
            data_re_out => mul_re_out(368),
            data_im_out => mul_im_out(368)
        );

 
    UMUL_369 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(369),
            data_im_in => first_stage_im_out(369),
            re_multiplicator => "1101010110011011", --- -0.662414550781 + j-0.749145507812
            im_multiplicator => "1101000000001110",
            data_re_out => mul_re_out(369),
            data_im_out => mul_im_out(369)
        );

 
    UMUL_370 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(370),
            data_im_in => first_stage_im_out(370),
            re_multiplicator => "1100111110001010", --- -0.757202148438 + j-0.653198242188
            im_multiplicator => "1101011000110010",
            data_re_out => mul_re_out(370),
            data_im_out => mul_im_out(370)
        );

 
    UMUL_371 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(371),
            data_im_in => first_stage_im_out(371),
            re_multiplicator => "1100101001011011", --- -0.838195800781 + j-0.545349121094
            im_multiplicator => "1101110100011001",
            data_re_out => mul_re_out(371),
            data_im_out => mul_im_out(371)
        );

 
    UMUL_372 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(372),
            data_im_in => first_stage_im_out(372),
            re_multiplicator => "1100011000100101", --- -0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(372),
            data_im_out => mul_im_out(372)
        );

 
    UMUL_373 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(373),
            data_im_in => first_stage_im_out(373),
            re_multiplicator => "1100001011111101", --- -0.953308105469 + j-0.302001953125
            im_multiplicator => "1110110010101100",
            data_re_out => mul_re_out(373),
            data_im_out => mul_im_out(373)
        );

 
    UMUL_374 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(374),
            data_im_in => first_stage_im_out(374),
            re_multiplicator => "1100000011110001", --- -0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(374),
            data_im_out => mul_im_out(374)
        );

 
    UMUL_375 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(375),
            data_im_in => first_stage_im_out(375),
            re_multiplicator => "1100000000001011", --- -0.999328613281 + j-0.0368041992188
            im_multiplicator => "1111110110100101",
            data_re_out => mul_re_out(375),
            data_im_out => mul_im_out(375)
        );

 
    UMUL_376 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(376),
            data_im_in => first_stage_im_out(376),
            re_multiplicator => "1100000001001111", --- -0.995178222656 + j0.0980224609375
            im_multiplicator => "0000011001000110",
            data_re_out => mul_re_out(376),
            data_im_out => mul_im_out(376)
        );

 
    UMUL_377 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(377),
            data_im_in => first_stage_im_out(377),
            re_multiplicator => "1100000110111011", --- -0.972961425781 + j0.231079101562
            im_multiplicator => "0000111011001010",
            data_re_out => mul_re_out(377),
            data_im_out => mul_im_out(377)
        );

 
    UMUL_378 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(378),
            data_im_in => first_stage_im_out(378),
            re_multiplicator => "1100010001001010", --- -0.932983398438 + j0.359924316406
            im_multiplicator => "0001011100001001",
            data_re_out => mul_re_out(378),
            data_im_out => mul_im_out(378)
        );

 
    UMUL_379 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(379),
            data_im_in => first_stage_im_out(379),
            re_multiplicator => "1100011111101110", --- -0.876098632812 + j0.482177734375
            im_multiplicator => "0001111011011100",
            data_re_out => mul_re_out(379),
            data_im_out => mul_im_out(379)
        );

 
    UMUL_380 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(380),
            data_im_in => first_stage_im_out(380),
            re_multiplicator => "1100110010011000", --- -0.80322265625 + j0.595703125
            im_multiplicator => "0010011000100000",
            data_re_out => mul_re_out(380),
            data_im_out => mul_im_out(380)
        );

 
    UMUL_381 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(381),
            data_im_in => first_stage_im_out(381),
            re_multiplicator => "1101001000110001", --- -0.715759277344 + j0.698364257812
            im_multiplicator => "0010110010110010",
            data_re_out => mul_re_out(381),
            data_im_out => mul_im_out(381)
        );

 
    UMUL_382 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(382),
            data_im_in => first_stage_im_out(382),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j0.788330078125
            im_multiplicator => "0011001001110100",
            data_re_out => mul_re_out(382),
            data_im_out => mul_im_out(382)
        );

 
    UMUL_383 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(383),
            data_im_in => first_stage_im_out(383),
            re_multiplicator => "1101111111000110", --- -0.503540039062 + j0.863952636719
            im_multiplicator => "0011011101001011",
            data_re_out => mul_re_out(383),
            data_im_out => mul_im_out(383)
        );

 
    UMUL_384 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(384),
            data_im_in => first_stage_im_out(384),
            data_re_out => mul_re_out(384),
            data_im_out => mul_im_out(384)
        );

 
    UMUL_385 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(385),
            data_im_in => first_stage_im_out(385),
            re_multiplicator => "0011111101001111", --- 0.989196777344 + j-0.146728515625
            im_multiplicator => "1111011010011100",
            data_re_out => mul_re_out(385),
            data_im_out => mul_im_out(385)
        );

 
    UMUL_386 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(386),
            data_im_in => first_stage_im_out(386),
            re_multiplicator => "0011110100111111", --- 0.956970214844 + j-0.290283203125
            im_multiplicator => "1110110101101100",
            data_re_out => mul_re_out(386),
            data_im_out => mul_im_out(386)
        );

 
    UMUL_387 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(387),
            data_im_in => first_stage_im_out(387),
            re_multiplicator => "0011100111011011", --- 0.903991699219 + j-0.427551269531
            im_multiplicator => "1110010010100011",
            data_re_out => mul_re_out(387),
            data_im_out => mul_im_out(387)
        );

 
    UMUL_388 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(388),
            data_im_in => first_stage_im_out(388),
            re_multiplicator => "0011010100110111", --- 0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(388),
            data_im_out => mul_im_out(388)
        );

 
    UMUL_389 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(389),
            data_im_in => first_stage_im_out(389),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(389),
            data_im_out => mul_im_out(389)
        );

 
    UMUL_390 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(390),
            data_im_in => first_stage_im_out(390),
            re_multiplicator => "0010100010011010", --- 0.634399414062 + j-0.773010253906
            im_multiplicator => "1100111010000111",
            data_re_out => mul_re_out(390),
            data_im_out => mul_im_out(390)
        );

 
    UMUL_391 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(391),
            data_im_in => first_stage_im_out(391),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(391),
            data_im_out => mul_im_out(391)
        );

 
    UMUL_392 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(392),
            data_im_in => first_stage_im_out(392),
            re_multiplicator => "0001100001111110", --- 0.382690429688 + j-0.923889160156
            im_multiplicator => "1100010011011111",
            data_re_out => mul_re_out(392),
            data_im_out => mul_im_out(392)
        );

 
    UMUL_393 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(393),
            data_im_in => first_stage_im_out(393),
            re_multiplicator => "0000111110001101", --- 0.242980957031 + j-0.970031738281
            im_multiplicator => "1100000111101011",
            data_re_out => mul_re_out(393),
            data_im_out => mul_im_out(393)
        );

 
    UMUL_394 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(394),
            data_im_in => first_stage_im_out(394),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(394),
            data_im_out => mul_im_out(394)
        );

 
    UMUL_395 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(395),
            data_im_in => first_stage_im_out(395),
            re_multiplicator => "1111110011011100", --- -0.049072265625 + j-0.998779296875
            im_multiplicator => "1100000000010100",
            data_re_out => mul_re_out(395),
            data_im_out => mul_im_out(395)
        );

 
    UMUL_396 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(396),
            data_im_in => first_stage_im_out(396),
            re_multiplicator => "1111001110000100", --- -0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(396),
            data_im_out => mul_im_out(396)
        );

 
    UMUL_397 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(397),
            data_im_in => first_stage_im_out(397),
            re_multiplicator => "1110101001110000", --- -0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(397),
            data_im_out => mul_im_out(397)
        );

 
    UMUL_398 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(398),
            data_im_in => first_stage_im_out(398),
            re_multiplicator => "1110000111010101", --- -0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(398),
            data_im_out => mul_im_out(398)
        );

 
    UMUL_399 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(399),
            data_im_in => first_stage_im_out(399),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(399),
            data_im_out => mul_im_out(399)
        );

 
    UMUL_400 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(400),
            data_im_in => first_stage_im_out(400),
            re_multiplicator => "1101001010111111", --- -0.707092285156 + j-0.707092285156
            im_multiplicator => "1101001010111111",
            data_re_out => mul_re_out(400),
            data_im_out => mul_im_out(400)
        );

 
    UMUL_401 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(401),
            data_im_in => first_stage_im_out(401),
            re_multiplicator => "1100110010011000", --- -0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(401),
            data_im_out => mul_im_out(401)
        );

 
    UMUL_402 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(402),
            data_im_in => first_stage_im_out(402),
            re_multiplicator => "1100011110001111", --- -0.881896972656 + j-0.471374511719
            im_multiplicator => "1110000111010101",
            data_re_out => mul_re_out(402),
            data_im_out => mul_im_out(402)
        );

 
    UMUL_403 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(403),
            data_im_in => first_stage_im_out(403),
            re_multiplicator => "1100001110111110", --- -0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(403),
            data_im_out => mul_im_out(403)
        );

 
    UMUL_404 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(404),
            data_im_in => first_stage_im_out(404),
            re_multiplicator => "1100000100111011", --- -0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(404),
            data_im_out => mul_im_out(404)
        );

 
    UMUL_405 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(405),
            data_im_in => first_stage_im_out(405),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(405),
            data_im_out => mul_im_out(405)
        );

 
    UMUL_406 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(406),
            data_im_in => first_stage_im_out(406),
            re_multiplicator => "1100000001001111", --- -0.995178222656 + j0.0980224609375
            im_multiplicator => "0000011001000110",
            data_re_out => mul_re_out(406),
            data_im_out => mul_im_out(406)
        );

 
    UMUL_407 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(407),
            data_im_in => first_stage_im_out(407),
            re_multiplicator => "1100000111101011", --- -0.970031738281 + j0.242980957031
            im_multiplicator => "0000111110001101",
            data_re_out => mul_re_out(407),
            data_im_out => mul_im_out(407)
        );

 
    UMUL_408 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(408),
            data_im_in => first_stage_im_out(408),
            re_multiplicator => "1100010011011111", --- -0.923889160156 + j0.382690429688
            im_multiplicator => "0001100001111110",
            data_re_out => mul_re_out(408),
            data_im_out => mul_im_out(408)
        );

 
    UMUL_409 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(409),
            data_im_in => first_stage_im_out(409),
            re_multiplicator => "1100100100011011", --- -0.857727050781 + j0.514099121094
            im_multiplicator => "0010000011100111",
            data_re_out => mul_re_out(409),
            data_im_out => mul_im_out(409)
        );

 
    UMUL_410 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(410),
            data_im_in => first_stage_im_out(410),
            re_multiplicator => "1100111010000111", --- -0.773010253906 + j0.634399414062
            im_multiplicator => "0010100010011010",
            data_re_out => mul_re_out(410),
            data_im_out => mul_im_out(410)
        );

 
    UMUL_411 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(411),
            data_im_in => first_stage_im_out(411),
            re_multiplicator => "1101010100000101", --- -0.671569824219 + j0.740966796875
            im_multiplicator => "0010111101101100",
            data_re_out => mul_re_out(411),
            data_im_out => mul_im_out(411)
        );

 
    UMUL_412 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(412),
            data_im_in => first_stage_im_out(412),
            re_multiplicator => "1101110001110010", --- -0.555541992188 + j0.831481933594
            im_multiplicator => "0011010100110111",
            data_re_out => mul_re_out(412),
            data_im_out => mul_im_out(412)
        );

 
    UMUL_413 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(413),
            data_im_in => first_stage_im_out(413),
            re_multiplicator => "1110010010100011", --- -0.427551269531 + j0.903991699219
            im_multiplicator => "0011100111011011",
            data_re_out => mul_re_out(413),
            data_im_out => mul_im_out(413)
        );

 
    UMUL_414 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(414),
            data_im_in => first_stage_im_out(414),
            re_multiplicator => "1110110101101100", --- -0.290283203125 + j0.956970214844
            im_multiplicator => "0011110100111111",
            data_re_out => mul_re_out(414),
            data_im_out => mul_im_out(414)
        );

 
    UMUL_415 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(415),
            data_im_in => first_stage_im_out(415),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j0.989196777344
            im_multiplicator => "0011111101001111",
            data_re_out => mul_re_out(415),
            data_im_out => mul_im_out(415)
        );

 
    UMUL_416 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(416),
            data_im_in => first_stage_im_out(416),
            data_re_out => mul_re_out(416),
            data_im_out => mul_im_out(416)
        );

 
    UMUL_417 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(417),
            data_im_in => first_stage_im_out(417),
            re_multiplicator => "0011111100110000", --- 0.9873046875 + j-0.158874511719
            im_multiplicator => "1111010111010101",
            data_re_out => mul_re_out(417),
            data_im_out => mul_im_out(417)
        );

 
    UMUL_418 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(418),
            data_im_in => first_stage_im_out(418),
            re_multiplicator => "0011110011000101", --- 0.949523925781 + j-0.313659667969
            im_multiplicator => "1110101111101101",
            data_re_out => mul_re_out(418),
            data_im_out => mul_im_out(418)
        );

 
    UMUL_419 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(419),
            data_im_in => first_stage_im_out(419),
            re_multiplicator => "0011100011001111", --- 0.887634277344 + j-0.460510253906
            im_multiplicator => "1110001010000111",
            data_re_out => mul_re_out(419),
            data_im_out => mul_im_out(419)
        );

 
    UMUL_420 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(420),
            data_im_in => first_stage_im_out(420),
            re_multiplicator => "0011001101101000", --- 0.80322265625 + j-0.595703125
            im_multiplicator => "1101100111100000",
            data_re_out => mul_re_out(420),
            data_im_out => mul_im_out(420)
        );

 
    UMUL_421 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(421),
            data_im_in => first_stage_im_out(421),
            re_multiplicator => "0010110010110010", --- 0.698364257812 + j-0.715759277344
            im_multiplicator => "1101001000110001",
            data_re_out => mul_re_out(421),
            data_im_out => mul_im_out(421)
        );

 
    UMUL_422 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(422),
            data_im_in => first_stage_im_out(422),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j-0.817565917969
            im_multiplicator => "1100101110101101",
            data_re_out => mul_re_out(422),
            data_im_out => mul_im_out(422)
        );

 
    UMUL_423 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(423),
            data_im_in => first_stage_im_out(423),
            re_multiplicator => "0001110000010010", --- 0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(423),
            data_im_out => mul_im_out(423)
        );

 
    UMUL_424 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(424),
            data_im_in => first_stage_im_out(424),
            re_multiplicator => "0001001010010100", --- 0.290283203125 + j-0.956970214844
            im_multiplicator => "1100001011000001",
            data_re_out => mul_re_out(424),
            data_im_out => mul_im_out(424)
        );

 
    UMUL_425 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(425),
            data_im_in => first_stage_im_out(425),
            re_multiplicator => "0000100010011101", --- 0.134582519531 + j-0.990905761719
            im_multiplicator => "1100000010010101",
            data_re_out => mul_re_out(425),
            data_im_out => mul_im_out(425)
        );

 
    UMUL_426 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(426),
            data_im_in => first_stage_im_out(426),
            re_multiplicator => "1111111001101110", --- -0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(426),
            data_im_out => mul_im_out(426)
        );

 
    UMUL_427 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(427),
            data_im_in => first_stage_im_out(427),
            re_multiplicator => "1111010001001001", --- -0.183044433594 + j-0.983093261719
            im_multiplicator => "1100000100010101",
            data_re_out => mul_re_out(427),
            data_im_out => mul_im_out(427)
        );

 
    UMUL_428 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(428),
            data_im_in => first_stage_im_out(428),
            re_multiplicator => "1110101001110000", --- -0.3369140625 + j-0.941528320312
            im_multiplicator => "1100001110111110",
            data_re_out => mul_re_out(428),
            data_im_out => mul_im_out(428)
        );

 
    UMUL_429 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(429),
            data_im_in => first_stage_im_out(429),
            re_multiplicator => "1110000100100100", --- -0.482177734375 + j-0.876098632812
            im_multiplicator => "1100011111101110",
            data_re_out => mul_re_out(429),
            data_im_out => mul_im_out(429)
        );

 
    UMUL_430 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(430),
            data_im_in => first_stage_im_out(430),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j-0.788330078125
            im_multiplicator => "1100110110001100",
            data_re_out => mul_re_out(430),
            data_im_out => mul_im_out(430)
        );

 
    UMUL_431 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(431),
            data_im_in => first_stage_im_out(431),
            re_multiplicator => "1101000100011100", --- -0.732666015625 + j-0.680603027344
            im_multiplicator => "1101010001110001",
            data_re_out => mul_re_out(431),
            data_im_out => mul_im_out(431)
        );

 
    UMUL_432 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(432),
            data_im_in => first_stage_im_out(432),
            re_multiplicator => "1100101011001001", --- -0.831481933594 + j-0.555541992188
            im_multiplicator => "1101110001110010",
            data_re_out => mul_re_out(432),
            data_im_out => mul_im_out(432)
        );

 
    UMUL_433 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(433),
            data_im_in => first_stage_im_out(433),
            re_multiplicator => "1100010111010000", --- -0.9091796875 + j-0.416442871094
            im_multiplicator => "1110010101011001",
            data_re_out => mul_re_out(433),
            data_im_out => mul_im_out(433)
        );

 
    UMUL_434 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(434),
            data_im_in => first_stage_im_out(434),
            re_multiplicator => "1100001001010001", --- -0.963806152344 + j-0.266723632812
            im_multiplicator => "1110111011101110",
            data_re_out => mul_re_out(434),
            data_im_out => mul_im_out(434)
        );

 
    UMUL_435 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(435),
            data_im_in => first_stage_im_out(435),
            re_multiplicator => "1100000001100100", --- -0.993896484375 + j-0.110229492188
            im_multiplicator => "1111100011110010",
            data_re_out => mul_re_out(435),
            data_im_out => mul_im_out(435)
        );

 
    UMUL_436 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(436),
            data_im_in => first_stage_im_out(436),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j0.049072265625
            im_multiplicator => "0000001100100100",
            data_re_out => mul_re_out(436),
            data_im_out => mul_im_out(436)
        );

 
    UMUL_437 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(437),
            data_im_in => first_stage_im_out(437),
            re_multiplicator => "1100000101100011", --- -0.978332519531 + j0.207092285156
            im_multiplicator => "0000110101000001",
            data_re_out => mul_re_out(437),
            data_im_out => mul_im_out(437)
        );

 
    UMUL_438 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(438),
            data_im_in => first_stage_im_out(438),
            re_multiplicator => "1100010001001010", --- -0.932983398438 + j0.359924316406
            im_multiplicator => "0001011100001001",
            data_re_out => mul_re_out(438),
            data_im_out => mul_im_out(438)
        );

 
    UMUL_439 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(439),
            data_im_in => first_stage_im_out(439),
            re_multiplicator => "1100100010110101", --- -0.863952636719 + j0.503540039062
            im_multiplicator => "0010000000111010",
            data_re_out => mul_re_out(439),
            data_im_out => mul_im_out(439)
        );

 
    UMUL_440 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(440),
            data_im_in => first_stage_im_out(440),
            re_multiplicator => "1100111010000111", --- -0.773010253906 + j0.634399414062
            im_multiplicator => "0010100010011010",
            data_re_out => mul_re_out(440),
            data_im_out => mul_im_out(440)
        );

 
    UMUL_441 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(441),
            data_im_in => first_stage_im_out(441),
            re_multiplicator => "1101010110011011", --- -0.662414550781 + j0.749145507812
            im_multiplicator => "0010111111110010",
            data_re_out => mul_re_out(441),
            data_im_out => mul_im_out(441)
        );

 
    UMUL_442 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(442),
            data_im_in => first_stage_im_out(442),
            re_multiplicator => "1101110111000011", --- -0.534973144531 + j0.844848632812
            im_multiplicator => "0011011000010010",
            data_re_out => mul_re_out(442),
            data_im_out => mul_im_out(442)
        );

 
    UMUL_443 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(443),
            data_im_in => first_stage_im_out(443),
            re_multiplicator => "1110011011001001", --- -0.393981933594 + j0.919128417969
            im_multiplicator => "0011101011010011",
            data_re_out => mul_re_out(443),
            data_im_out => mul_im_out(443)
        );

 
    UMUL_444 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(444),
            data_im_in => first_stage_im_out(444),
            re_multiplicator => "1111000001110011", --- -0.242980957031 + j0.970031738281
            im_multiplicator => "0011111000010101",
            data_re_out => mul_re_out(444),
            data_im_out => mul_im_out(444)
        );

 
    UMUL_445 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(445),
            data_im_in => first_stage_im_out(445),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j0.996337890625
            im_multiplicator => "0011111111000100",
            data_re_out => mul_re_out(445),
            data_im_out => mul_im_out(445)
        );

 
    UMUL_446 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(446),
            data_im_in => first_stage_im_out(446),
            re_multiplicator => "0000010010110101", --- 0.0735473632812 + j0.997314453125
            im_multiplicator => "0011111111010100",
            data_re_out => mul_re_out(446),
            data_im_out => mul_im_out(446)
        );

 
    UMUL_447 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(447),
            data_im_in => first_stage_im_out(447),
            re_multiplicator => "0000111011001010", --- 0.231079101562 + j0.972961425781
            im_multiplicator => "0011111001000101",
            data_re_out => mul_re_out(447),
            data_im_out => mul_im_out(447)
        );

 
    UMUL_448 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(448),
            data_im_in => first_stage_im_out(448),
            data_re_out => mul_re_out(448),
            data_im_out => mul_im_out(448)
        );

 
    UMUL_449 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(449),
            data_im_in => first_stage_im_out(449),
            re_multiplicator => "0011111100001111", --- 0.985290527344 + j-0.170959472656
            im_multiplicator => "1111010100001111",
            data_re_out => mul_re_out(449),
            data_im_out => mul_im_out(449)
        );

 
    UMUL_450 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(450),
            data_im_in => first_stage_im_out(450),
            re_multiplicator => "0011110001000010", --- 0.941528320312 + j-0.3369140625
            im_multiplicator => "1110101001110000",
            data_re_out => mul_re_out(450),
            data_im_out => mul_im_out(450)
        );

 
    UMUL_451 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(451),
            data_im_in => first_stage_im_out(451),
            re_multiplicator => "0011011110110000", --- 0.8701171875 + j-0.492919921875
            im_multiplicator => "1110000001110100",
            data_re_out => mul_re_out(451),
            data_im_out => mul_im_out(451)
        );

 
    UMUL_452 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(452),
            data_im_in => first_stage_im_out(452),
            re_multiplicator => "0011000101111001", --- 0.773010253906 + j-0.634399414062
            im_multiplicator => "1101011101100110",
            data_re_out => mul_re_out(452),
            data_im_out => mul_im_out(452)
        );

 
    UMUL_453 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(453),
            data_im_in => first_stage_im_out(453),
            re_multiplicator => "0010100111001110", --- 0.653198242188 + j-0.757202148438
            im_multiplicator => "1100111110001010",
            data_re_out => mul_re_out(453),
            data_im_out => mul_im_out(453)
        );

 
    UMUL_454 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(454),
            data_im_in => first_stage_im_out(454),
            re_multiplicator => "0010000011100111", --- 0.514099121094 + j-0.857727050781
            im_multiplicator => "1100100100011011",
            data_re_out => mul_re_out(454),
            data_im_out => mul_im_out(454)
        );

 
    UMUL_455 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(455),
            data_im_in => first_stage_im_out(455),
            re_multiplicator => "0001011100001001", --- 0.359924316406 + j-0.932983398438
            im_multiplicator => "1100010001001010",
            data_re_out => mul_re_out(455),
            data_im_out => mul_im_out(455)
        );

 
    UMUL_456 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(456),
            data_im_in => first_stage_im_out(456),
            re_multiplicator => "0000110001111100", --- 0.195068359375 + j-0.980773925781
            im_multiplicator => "1100000100111011",
            data_re_out => mul_re_out(456),
            data_im_out => mul_im_out(456)
        );

 
    UMUL_457 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(457),
            data_im_in => first_stage_im_out(457),
            re_multiplicator => "0000000110010010", --- 0.0245361328125 + j-0.999694824219
            im_multiplicator => "1100000000000101",
            data_re_out => mul_re_out(457),
            data_im_out => mul_im_out(457)
        );

 
    UMUL_458 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(458),
            data_im_in => first_stage_im_out(458),
            re_multiplicator => "1111011010011100", --- -0.146728515625 + j-0.989196777344
            im_multiplicator => "1100000010110001",
            data_re_out => mul_re_out(458),
            data_im_out => mul_im_out(458)
        );

 
    UMUL_459 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(459),
            data_im_in => first_stage_im_out(459),
            re_multiplicator => "1110101111101101", --- -0.313659667969 + j-0.949523925781
            im_multiplicator => "1100001100111011",
            data_re_out => mul_re_out(459),
            data_im_out => mul_im_out(459)
        );

 
    UMUL_460 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(460),
            data_im_in => first_stage_im_out(460),
            re_multiplicator => "1110000111010101", --- -0.471374511719 + j-0.881896972656
            im_multiplicator => "1100011110001111",
            data_re_out => mul_re_out(460),
            data_im_out => mul_im_out(460)
        );

 
    UMUL_461 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(461),
            data_im_in => first_stage_im_out(461),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j-0.788330078125
            im_multiplicator => "1100110110001100",
            data_re_out => mul_re_out(461),
            data_im_out => mul_im_out(461)
        );

 
    UMUL_462 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(462),
            data_im_in => first_stage_im_out(462),
            re_multiplicator => "1101000010010100", --- -0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(462),
            data_im_out => mul_im_out(462)
        );

 
    UMUL_463 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(463),
            data_im_in => first_stage_im_out(463),
            re_multiplicator => "1100100111101110", --- -0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(463),
            data_im_out => mul_im_out(463)
        );

 
    UMUL_464 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(464),
            data_im_in => first_stage_im_out(464),
            re_multiplicator => "1100010011011111", --- -0.923889160156 + j-0.382690429688
            im_multiplicator => "1110011110000010",
            data_re_out => mul_re_out(464),
            data_im_out => mul_im_out(464)
        );

 
    UMUL_465 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(465),
            data_im_in => first_stage_im_out(465),
            re_multiplicator => "1100000110001110", --- -0.975708007812 + j-0.219116210938
            im_multiplicator => "1111000111111010",
            data_re_out => mul_re_out(465),
            data_im_out => mul_im_out(465)
        );

 
    UMUL_466 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(466),
            data_im_in => first_stage_im_out(466),
            re_multiplicator => "1100000000010100", --- -0.998779296875 + j-0.049072265625
            im_multiplicator => "1111110011011100",
            data_re_out => mul_re_out(466),
            data_im_out => mul_im_out(466)
        );

 
    UMUL_467 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(467),
            data_im_in => first_stage_im_out(467),
            re_multiplicator => "1100000001111011", --- -0.992492675781 + j0.122436523438
            im_multiplicator => "0000011111010110",
            data_re_out => mul_re_out(467),
            data_im_out => mul_im_out(467)
        );

 
    UMUL_468 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(468),
            data_im_in => first_stage_im_out(468),
            re_multiplicator => "1100001011000001", --- -0.956970214844 + j0.290283203125
            im_multiplicator => "0001001010010100",
            data_re_out => mul_re_out(468),
            data_im_out => mul_im_out(468)
        );

 
    UMUL_469 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(469),
            data_im_in => first_stage_im_out(469),
            re_multiplicator => "1100011011010101", --- -0.893249511719 + j0.449584960938
            im_multiplicator => "0001110011000110",
            data_re_out => mul_re_out(469),
            data_im_out => mul_im_out(469)
        );

 
    UMUL_470 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(470),
            data_im_in => first_stage_im_out(470),
            re_multiplicator => "1100110010011000", --- -0.80322265625 + j0.595703125
            im_multiplicator => "0010011000100000",
            data_re_out => mul_re_out(470),
            data_im_out => mul_im_out(470)
        );

 
    UMUL_471 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(471),
            data_im_in => first_stage_im_out(471),
            re_multiplicator => "1101001111011111", --- -0.689514160156 + j0.724243164062
            im_multiplicator => "0010111001011010",
            data_re_out => mul_re_out(471),
            data_im_out => mul_im_out(471)
        );

 
    UMUL_472 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(472),
            data_im_in => first_stage_im_out(472),
            re_multiplicator => "1101110001110010", --- -0.555541992188 + j0.831481933594
            im_multiplicator => "0011010100110111",
            data_re_out => mul_re_out(472),
            data_im_out => mul_im_out(472)
        );

 
    UMUL_473 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(473),
            data_im_in => first_stage_im_out(473),
            re_multiplicator => "1110011000010001", --- -0.405212402344 + j0.914184570312
            im_multiplicator => "0011101010000010",
            data_re_out => mul_re_out(473),
            data_im_out => mul_im_out(473)
        );

 
    UMUL_474 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(474),
            data_im_in => first_stage_im_out(474),
            re_multiplicator => "1111000001110011", --- -0.242980957031 + j0.970031738281
            im_multiplicator => "0011111000010101",
            data_re_out => mul_re_out(474),
            data_im_out => mul_im_out(474)
        );

 
    UMUL_475 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(475),
            data_im_in => first_stage_im_out(475),
            re_multiplicator => "1111101101001011", --- -0.0735473632812 + j0.997314453125
            im_multiplicator => "0011111111010100",
            data_re_out => mul_re_out(475),
            data_im_out => mul_im_out(475)
        );

 
    UMUL_476 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(476),
            data_im_in => first_stage_im_out(476),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j0.995178222656
            im_multiplicator => "0011111110110001",
            data_re_out => mul_re_out(476),
            data_im_out => mul_im_out(476)
        );

 
    UMUL_477 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(477),
            data_im_in => first_stage_im_out(477),
            re_multiplicator => "0001000100010010", --- 0.266723632812 + j0.963806152344
            im_multiplicator => "0011110110101111",
            data_re_out => mul_re_out(477),
            data_im_out => mul_im_out(477)
        );

 
    UMUL_478 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(478),
            data_im_in => first_stage_im_out(478),
            re_multiplicator => "0001101101011101", --- 0.427551269531 + j0.903991699219
            im_multiplicator => "0011100111011011",
            data_re_out => mul_re_out(478),
            data_im_out => mul_im_out(478)
        );

 
    UMUL_479 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(479),
            data_im_in => first_stage_im_out(479),
            re_multiplicator => "0010010011011010", --- 0.575805664062 + j0.817565917969
            im_multiplicator => "0011010001010011",
            data_re_out => mul_re_out(479),
            data_im_out => mul_im_out(479)
        );

 
    UMUL_480 : multiplier_mul1
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(480),
            data_im_in => first_stage_im_out(480),
            data_re_out => mul_re_out(480),
            data_im_out => mul_im_out(480)
        );

 
    UMUL_481 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(481),
            data_im_in => first_stage_im_out(481),
            re_multiplicator => "0011111011101011", --- 0.983093261719 + j-0.183044433594
            im_multiplicator => "1111010001001001",
            data_re_out => mul_re_out(481),
            data_im_out => mul_im_out(481)
        );

 
    UMUL_482 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(482),
            data_im_in => first_stage_im_out(482),
            re_multiplicator => "0011101110110110", --- 0.932983398438 + j-0.359924316406
            im_multiplicator => "1110100011110111",
            data_re_out => mul_re_out(482),
            data_im_out => mul_im_out(482)
        );

 
    UMUL_483 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(483),
            data_im_in => first_stage_im_out(483),
            re_multiplicator => "0011011001111101", --- 0.851379394531 + j-0.524597167969
            im_multiplicator => "1101111001101101",
            data_re_out => mul_re_out(483),
            data_im_out => mul_im_out(483)
        );

 
    UMUL_484 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(484),
            data_im_in => first_stage_im_out(484),
            re_multiplicator => "0010111101101100", --- 0.740966796875 + j-0.671569824219
            im_multiplicator => "1101010100000101",
            data_re_out => mul_re_out(484),
            data_im_out => mul_im_out(484)
        );

 
    UMUL_485 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(485),
            data_im_in => first_stage_im_out(485),
            re_multiplicator => "0010011011000001", --- 0.605529785156 + j-0.795837402344
            im_multiplicator => "1100110100010001",
            data_re_out => mul_re_out(485),
            data_im_out => mul_im_out(485)
        );

 
    UMUL_486 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(486),
            data_im_in => first_stage_im_out(486),
            re_multiplicator => "0001110011000110", --- 0.449584960938 + j-0.893249511719
            im_multiplicator => "1100011011010101",
            data_re_out => mul_re_out(486),
            data_im_out => mul_im_out(486)
        );

 
    UMUL_487 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(487),
            data_im_in => first_stage_im_out(487),
            re_multiplicator => "0001000111010011", --- 0.278503417969 + j-0.96044921875
            im_multiplicator => "1100001010001000",
            data_re_out => mul_re_out(487),
            data_im_out => mul_im_out(487)
        );

 
    UMUL_488 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(488),
            data_im_in => first_stage_im_out(488),
            re_multiplicator => "0000011001000110", --- 0.0980224609375 + j-0.995178222656
            im_multiplicator => "1100000001001111",
            data_re_out => mul_re_out(488),
            data_im_out => mul_im_out(488)
        );

 
    UMUL_489 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(489),
            data_im_in => first_stage_im_out(489),
            re_multiplicator => "1111101010000010", --- -0.0858154296875 + j-0.996337890625
            im_multiplicator => "1100000000111100",
            data_re_out => mul_re_out(489),
            data_im_out => mul_im_out(489)
        );

 
    UMUL_490 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(490),
            data_im_in => first_stage_im_out(490),
            re_multiplicator => "1110111011101110", --- -0.266723632812 + j-0.963806152344
            im_multiplicator => "1100001001010001",
            data_re_out => mul_re_out(490),
            data_im_out => mul_im_out(490)
        );

 
    UMUL_491 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(491),
            data_im_in => first_stage_im_out(491),
            re_multiplicator => "1110001111101110", --- -0.438598632812 + j-0.898681640625
            im_multiplicator => "1100011001111100",
            data_re_out => mul_re_out(491),
            data_im_out => mul_im_out(491)
        );

 
    UMUL_492 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(492),
            data_im_in => first_stage_im_out(492),
            re_multiplicator => "1101100111100000", --- -0.595703125 + j-0.80322265625
            im_multiplicator => "1100110010011000",
            data_re_out => mul_re_out(492),
            data_im_out => mul_im_out(492)
        );

 
    UMUL_493 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(493),
            data_im_in => first_stage_im_out(493),
            re_multiplicator => "1101000100011100", --- -0.732666015625 + j-0.680603027344
            im_multiplicator => "1101010001110001",
            data_re_out => mul_re_out(493),
            data_im_out => mul_im_out(493)
        );

 
    UMUL_494 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(494),
            data_im_in => first_stage_im_out(494),
            re_multiplicator => "1100100111101110", --- -0.844848632812 + j-0.534973144531
            im_multiplicator => "1101110111000011",
            data_re_out => mul_re_out(494),
            data_im_out => mul_im_out(494)
        );

 
    UMUL_495 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(495),
            data_im_in => first_stage_im_out(495),
            re_multiplicator => "1100010010010011", --- -0.928527832031 + j-0.371337890625
            im_multiplicator => "1110100000111100",
            data_re_out => mul_re_out(495),
            data_im_out => mul_im_out(495)
        );

 
    UMUL_496 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(496),
            data_im_in => first_stage_im_out(496),
            re_multiplicator => "1100000100111011", --- -0.980773925781 + j-0.195068359375
            im_multiplicator => "1111001110000100",
            data_re_out => mul_re_out(496),
            data_im_out => mul_im_out(496)
        );

 
    UMUL_497 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(497),
            data_im_in => first_stage_im_out(497),
            re_multiplicator => "1100000000000001", --- -0.999938964844 + j-0.0122680664062
            im_multiplicator => "1111111100110111",
            data_re_out => mul_re_out(497),
            data_im_out => mul_im_out(497)
        );

 
    UMUL_498 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(498),
            data_im_in => first_stage_im_out(498),
            re_multiplicator => "1100000011110001", --- -0.985290527344 + j0.170959472656
            im_multiplicator => "0000101011110001",
            data_re_out => mul_re_out(498),
            data_im_out => mul_im_out(498)
        );

 
    UMUL_499 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(499),
            data_im_in => first_stage_im_out(499),
            re_multiplicator => "1100010000000011", --- -0.937316894531 + j0.348388671875
            im_multiplicator => "0001011001001100",
            data_re_out => mul_re_out(499),
            data_im_out => mul_im_out(499)
        );

 
    UMUL_500 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(500),
            data_im_in => first_stage_im_out(500),
            re_multiplicator => "1100100100011011", --- -0.857727050781 + j0.514099121094
            im_multiplicator => "0010000011100111",
            data_re_out => mul_re_out(500),
            data_im_out => mul_im_out(500)
        );

 
    UMUL_501 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(501),
            data_im_in => first_stage_im_out(501),
            re_multiplicator => "1101000000001110", --- -0.749145507812 + j0.662414550781
            im_multiplicator => "0010101001100101",
            data_re_out => mul_re_out(501),
            data_im_out => mul_im_out(501)
        );

 
    UMUL_502 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(502),
            data_im_in => first_stage_im_out(502),
            re_multiplicator => "1101100010100000", --- -0.615234375 + j0.788330078125
            im_multiplicator => "0011001001110100",
            data_re_out => mul_re_out(502),
            data_im_out => mul_im_out(502)
        );

 
    UMUL_503 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(503),
            data_im_in => first_stage_im_out(503),
            re_multiplicator => "1110001010000111", --- -0.460510253906 + j0.887634277344
            im_multiplicator => "0011100011001111",
            data_re_out => mul_re_out(503),
            data_im_out => mul_im_out(503)
        );

 
    UMUL_504 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(504),
            data_im_in => first_stage_im_out(504),
            re_multiplicator => "1110110101101100", --- -0.290283203125 + j0.956970214844
            im_multiplicator => "0011110100111111",
            data_re_out => mul_re_out(504),
            data_im_out => mul_im_out(504)
        );

 
    UMUL_505 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(505),
            data_im_in => first_stage_im_out(505),
            re_multiplicator => "1111100011110010", --- -0.110229492188 + j0.993896484375
            im_multiplicator => "0011111110011100",
            data_re_out => mul_re_out(505),
            data_im_out => mul_im_out(505)
        );

 
    UMUL_506 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(506),
            data_im_in => first_stage_im_out(506),
            re_multiplicator => "0000010010110101", --- 0.0735473632812 + j0.997314453125
            im_multiplicator => "0011111111010100",
            data_re_out => mul_re_out(506),
            data_im_out => mul_im_out(506)
        );

 
    UMUL_507 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(507),
            data_im_in => first_stage_im_out(507),
            re_multiplicator => "0001000001010000", --- 0.2548828125 + j0.966979980469
            im_multiplicator => "0011110111100011",
            data_re_out => mul_re_out(507),
            data_im_out => mul_im_out(507)
        );

 
    UMUL_508 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(508),
            data_im_in => first_stage_im_out(508),
            re_multiplicator => "0001101101011101", --- 0.427551269531 + j0.903991699219
            im_multiplicator => "0011100111011011",
            data_re_out => mul_re_out(508),
            data_im_out => mul_im_out(508)
        );

 
    UMUL_509 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(509),
            data_im_in => first_stage_im_out(509),
            re_multiplicator => "0010010101111110", --- 0.585815429688 + j0.810485839844
            im_multiplicator => "0011001111011111",
            data_re_out => mul_re_out(509),
            data_im_out => mul_im_out(509)
        );

 
    UMUL_510 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(510),
            data_im_in => first_stage_im_out(510),
            re_multiplicator => "0010111001011010", --- 0.724243164062 + j0.689514160156
            im_multiplicator => "0010110000100001",
            data_re_out => mul_re_out(510),
            data_im_out => mul_im_out(510)
        );

 
    UMUL_511 : complex_multiplier
    generic map(
            ctrl_start => (ctrl_start+4) mod 16
        )
    port map(
            clk => clk,
            rst => rst,
            ce => ce,
            bypass => bypass(5),
            ctrl_delay => ctrl_delay,
            data_re_in => first_stage_re_out(511),
            data_im_in => first_stage_im_out(511),
            re_multiplicator => "0011010110100101", --- 0.838195800781 + j0.545349121094
            im_multiplicator => "0010001011100111",
            data_re_out => mul_re_out(511),
            data_im_out => mul_im_out(511)
        );

end Behavioral;
