library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity fft_pt2048 is
    PORT (
        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        ctrl           : IN STD_LOGIC;

        data_re_in:in std_logic_vector(2047 downto 0);
        data_im_in:in std_logic_vector(2047 downto 0);

        data_re_out:out std_logic_vector(2047 downto 0);
        data_im_out:out std_logic_vector(2047 downto 0)
    );
end fft_pt2048;

architecture Behavioral of fft_pt2048 is

component fft_pt32 is
    PORT (
        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        ctrl           : IN STD_LOGIC;

        data_re_in:in std_logic_vector(31 downto 0);
        data_im_in:in std_logic_vector(31 downto 0);

        data_re_out:out std_logic_vector(31 downto 0);
        data_im_out:out std_logic_vector(31 downto 0)
    );
end component;

component fft_pt64 is
    PORT (
        clk            : IN STD_LOGIC;
        rst            : IN STD_LOGIC;
        ce             : IN STD_LOGIC;
        ctrl           : IN STD_LOGIC;

        data_re_in     : in std_logic_vector(63 downto 0);
        data_im_in     : in std_logic_vector(63 downto 0);

        data_re_out     : out std_logic_vector(63 downto 0);
        data_im_out     : out std_logic_vector(63 downto 0)
    );
end component;

component complex_multiplier is
    GENERIC (
        re_multiplicator : INTEGER;
        im_multiplicator : INTEGER
    );
    PORT (
        clk             : IN std_logic;
        rst             : IN std_logic;
        ce              : IN std_logic;
        ctrl            : IN STD_LOGIC;
        data_re_in      : IN std_logic;
        data_im_in      : IN std_logic;
        product_re_out  : OUT STD_LOGIC;
        product_im_out  : OUT STD_LOGIC
    );
end component;

component Dff_regN is
    GENERIC( N: INTEGER );
    Port ( D : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           ce  : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           Q : out  STD_LOGIC);
end component;

component shifter is
    port(
            clk            : IN STD_LOGIC;
            rst            : IN STD_LOGIC;
            ce             : IN STD_LOGIC;
            ctrl           : IN STD_LOGIC;
            data_in:in std_logic;
            data_out:out std_logic
        );
end component;

signal first_stage_re_out, first_stage_im_out: std_logic_vector(2047 downto 0);
signal mul_re_out, mul_im_out : std_logic_vector(2047 downto 0);
signal shifter_re,shifter_im:std_logic_vector(2047 downto 0);
SIGNAL ctrl_delay : std_logic;

begin
    UDELAY_CTRL : Dff_regN
    generic map(N=>3)
    port map(
            D=>ctrl,
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>ctrl_delay
        );

    --- left-hand-side processors
    ULFFT_PT32_0 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(0),
            data_re_in(1)=>data_re_in(64),
            data_re_in(2)=>data_re_in(128),
            data_re_in(3)=>data_re_in(192),
            data_re_in(4)=>data_re_in(256),
            data_re_in(5)=>data_re_in(320),
            data_re_in(6)=>data_re_in(384),
            data_re_in(7)=>data_re_in(448),
            data_re_in(8)=>data_re_in(512),
            data_re_in(9)=>data_re_in(576),
            data_re_in(10)=>data_re_in(640),
            data_re_in(11)=>data_re_in(704),
            data_re_in(12)=>data_re_in(768),
            data_re_in(13)=>data_re_in(832),
            data_re_in(14)=>data_re_in(896),
            data_re_in(15)=>data_re_in(960),
            data_re_in(16)=>data_re_in(1024),
            data_re_in(17)=>data_re_in(1088),
            data_re_in(18)=>data_re_in(1152),
            data_re_in(19)=>data_re_in(1216),
            data_re_in(20)=>data_re_in(1280),
            data_re_in(21)=>data_re_in(1344),
            data_re_in(22)=>data_re_in(1408),
            data_re_in(23)=>data_re_in(1472),
            data_re_in(24)=>data_re_in(1536),
            data_re_in(25)=>data_re_in(1600),
            data_re_in(26)=>data_re_in(1664),
            data_re_in(27)=>data_re_in(1728),
            data_re_in(28)=>data_re_in(1792),
            data_re_in(29)=>data_re_in(1856),
            data_re_in(30)=>data_re_in(1920),
            data_re_in(31)=>data_re_in(1984),
            data_im_in(0)=>data_im_in(0),
            data_im_in(1)=>data_im_in(64),
            data_im_in(2)=>data_im_in(128),
            data_im_in(3)=>data_im_in(192),
            data_im_in(4)=>data_im_in(256),
            data_im_in(5)=>data_im_in(320),
            data_im_in(6)=>data_im_in(384),
            data_im_in(7)=>data_im_in(448),
            data_im_in(8)=>data_im_in(512),
            data_im_in(9)=>data_im_in(576),
            data_im_in(10)=>data_im_in(640),
            data_im_in(11)=>data_im_in(704),
            data_im_in(12)=>data_im_in(768),
            data_im_in(13)=>data_im_in(832),
            data_im_in(14)=>data_im_in(896),
            data_im_in(15)=>data_im_in(960),
            data_im_in(16)=>data_im_in(1024),
            data_im_in(17)=>data_im_in(1088),
            data_im_in(18)=>data_im_in(1152),
            data_im_in(19)=>data_im_in(1216),
            data_im_in(20)=>data_im_in(1280),
            data_im_in(21)=>data_im_in(1344),
            data_im_in(22)=>data_im_in(1408),
            data_im_in(23)=>data_im_in(1472),
            data_im_in(24)=>data_im_in(1536),
            data_im_in(25)=>data_im_in(1600),
            data_im_in(26)=>data_im_in(1664),
            data_im_in(27)=>data_im_in(1728),
            data_im_in(28)=>data_im_in(1792),
            data_im_in(29)=>data_im_in(1856),
            data_im_in(30)=>data_im_in(1920),
            data_im_in(31)=>data_im_in(1984),
            data_re_out=>first_stage_re_out(31 downto 0),
            data_im_out=>first_stage_im_out(31 downto 0)
        );

    ULFFT_PT32_1 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(1),
            data_re_in(1)=>data_re_in(65),
            data_re_in(2)=>data_re_in(129),
            data_re_in(3)=>data_re_in(193),
            data_re_in(4)=>data_re_in(257),
            data_re_in(5)=>data_re_in(321),
            data_re_in(6)=>data_re_in(385),
            data_re_in(7)=>data_re_in(449),
            data_re_in(8)=>data_re_in(513),
            data_re_in(9)=>data_re_in(577),
            data_re_in(10)=>data_re_in(641),
            data_re_in(11)=>data_re_in(705),
            data_re_in(12)=>data_re_in(769),
            data_re_in(13)=>data_re_in(833),
            data_re_in(14)=>data_re_in(897),
            data_re_in(15)=>data_re_in(961),
            data_re_in(16)=>data_re_in(1025),
            data_re_in(17)=>data_re_in(1089),
            data_re_in(18)=>data_re_in(1153),
            data_re_in(19)=>data_re_in(1217),
            data_re_in(20)=>data_re_in(1281),
            data_re_in(21)=>data_re_in(1345),
            data_re_in(22)=>data_re_in(1409),
            data_re_in(23)=>data_re_in(1473),
            data_re_in(24)=>data_re_in(1537),
            data_re_in(25)=>data_re_in(1601),
            data_re_in(26)=>data_re_in(1665),
            data_re_in(27)=>data_re_in(1729),
            data_re_in(28)=>data_re_in(1793),
            data_re_in(29)=>data_re_in(1857),
            data_re_in(30)=>data_re_in(1921),
            data_re_in(31)=>data_re_in(1985),
            data_im_in(0)=>data_im_in(1),
            data_im_in(1)=>data_im_in(65),
            data_im_in(2)=>data_im_in(129),
            data_im_in(3)=>data_im_in(193),
            data_im_in(4)=>data_im_in(257),
            data_im_in(5)=>data_im_in(321),
            data_im_in(6)=>data_im_in(385),
            data_im_in(7)=>data_im_in(449),
            data_im_in(8)=>data_im_in(513),
            data_im_in(9)=>data_im_in(577),
            data_im_in(10)=>data_im_in(641),
            data_im_in(11)=>data_im_in(705),
            data_im_in(12)=>data_im_in(769),
            data_im_in(13)=>data_im_in(833),
            data_im_in(14)=>data_im_in(897),
            data_im_in(15)=>data_im_in(961),
            data_im_in(16)=>data_im_in(1025),
            data_im_in(17)=>data_im_in(1089),
            data_im_in(18)=>data_im_in(1153),
            data_im_in(19)=>data_im_in(1217),
            data_im_in(20)=>data_im_in(1281),
            data_im_in(21)=>data_im_in(1345),
            data_im_in(22)=>data_im_in(1409),
            data_im_in(23)=>data_im_in(1473),
            data_im_in(24)=>data_im_in(1537),
            data_im_in(25)=>data_im_in(1601),
            data_im_in(26)=>data_im_in(1665),
            data_im_in(27)=>data_im_in(1729),
            data_im_in(28)=>data_im_in(1793),
            data_im_in(29)=>data_im_in(1857),
            data_im_in(30)=>data_im_in(1921),
            data_im_in(31)=>data_im_in(1985),
            data_re_out=>first_stage_re_out(63 downto 32),
            data_im_out=>first_stage_im_out(63 downto 32)
        );

    ULFFT_PT32_2 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(2),
            data_re_in(1)=>data_re_in(66),
            data_re_in(2)=>data_re_in(130),
            data_re_in(3)=>data_re_in(194),
            data_re_in(4)=>data_re_in(258),
            data_re_in(5)=>data_re_in(322),
            data_re_in(6)=>data_re_in(386),
            data_re_in(7)=>data_re_in(450),
            data_re_in(8)=>data_re_in(514),
            data_re_in(9)=>data_re_in(578),
            data_re_in(10)=>data_re_in(642),
            data_re_in(11)=>data_re_in(706),
            data_re_in(12)=>data_re_in(770),
            data_re_in(13)=>data_re_in(834),
            data_re_in(14)=>data_re_in(898),
            data_re_in(15)=>data_re_in(962),
            data_re_in(16)=>data_re_in(1026),
            data_re_in(17)=>data_re_in(1090),
            data_re_in(18)=>data_re_in(1154),
            data_re_in(19)=>data_re_in(1218),
            data_re_in(20)=>data_re_in(1282),
            data_re_in(21)=>data_re_in(1346),
            data_re_in(22)=>data_re_in(1410),
            data_re_in(23)=>data_re_in(1474),
            data_re_in(24)=>data_re_in(1538),
            data_re_in(25)=>data_re_in(1602),
            data_re_in(26)=>data_re_in(1666),
            data_re_in(27)=>data_re_in(1730),
            data_re_in(28)=>data_re_in(1794),
            data_re_in(29)=>data_re_in(1858),
            data_re_in(30)=>data_re_in(1922),
            data_re_in(31)=>data_re_in(1986),
            data_im_in(0)=>data_im_in(2),
            data_im_in(1)=>data_im_in(66),
            data_im_in(2)=>data_im_in(130),
            data_im_in(3)=>data_im_in(194),
            data_im_in(4)=>data_im_in(258),
            data_im_in(5)=>data_im_in(322),
            data_im_in(6)=>data_im_in(386),
            data_im_in(7)=>data_im_in(450),
            data_im_in(8)=>data_im_in(514),
            data_im_in(9)=>data_im_in(578),
            data_im_in(10)=>data_im_in(642),
            data_im_in(11)=>data_im_in(706),
            data_im_in(12)=>data_im_in(770),
            data_im_in(13)=>data_im_in(834),
            data_im_in(14)=>data_im_in(898),
            data_im_in(15)=>data_im_in(962),
            data_im_in(16)=>data_im_in(1026),
            data_im_in(17)=>data_im_in(1090),
            data_im_in(18)=>data_im_in(1154),
            data_im_in(19)=>data_im_in(1218),
            data_im_in(20)=>data_im_in(1282),
            data_im_in(21)=>data_im_in(1346),
            data_im_in(22)=>data_im_in(1410),
            data_im_in(23)=>data_im_in(1474),
            data_im_in(24)=>data_im_in(1538),
            data_im_in(25)=>data_im_in(1602),
            data_im_in(26)=>data_im_in(1666),
            data_im_in(27)=>data_im_in(1730),
            data_im_in(28)=>data_im_in(1794),
            data_im_in(29)=>data_im_in(1858),
            data_im_in(30)=>data_im_in(1922),
            data_im_in(31)=>data_im_in(1986),
            data_re_out=>first_stage_re_out(95 downto 64),
            data_im_out=>first_stage_im_out(95 downto 64)
        );

    ULFFT_PT32_3 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(3),
            data_re_in(1)=>data_re_in(67),
            data_re_in(2)=>data_re_in(131),
            data_re_in(3)=>data_re_in(195),
            data_re_in(4)=>data_re_in(259),
            data_re_in(5)=>data_re_in(323),
            data_re_in(6)=>data_re_in(387),
            data_re_in(7)=>data_re_in(451),
            data_re_in(8)=>data_re_in(515),
            data_re_in(9)=>data_re_in(579),
            data_re_in(10)=>data_re_in(643),
            data_re_in(11)=>data_re_in(707),
            data_re_in(12)=>data_re_in(771),
            data_re_in(13)=>data_re_in(835),
            data_re_in(14)=>data_re_in(899),
            data_re_in(15)=>data_re_in(963),
            data_re_in(16)=>data_re_in(1027),
            data_re_in(17)=>data_re_in(1091),
            data_re_in(18)=>data_re_in(1155),
            data_re_in(19)=>data_re_in(1219),
            data_re_in(20)=>data_re_in(1283),
            data_re_in(21)=>data_re_in(1347),
            data_re_in(22)=>data_re_in(1411),
            data_re_in(23)=>data_re_in(1475),
            data_re_in(24)=>data_re_in(1539),
            data_re_in(25)=>data_re_in(1603),
            data_re_in(26)=>data_re_in(1667),
            data_re_in(27)=>data_re_in(1731),
            data_re_in(28)=>data_re_in(1795),
            data_re_in(29)=>data_re_in(1859),
            data_re_in(30)=>data_re_in(1923),
            data_re_in(31)=>data_re_in(1987),
            data_im_in(0)=>data_im_in(3),
            data_im_in(1)=>data_im_in(67),
            data_im_in(2)=>data_im_in(131),
            data_im_in(3)=>data_im_in(195),
            data_im_in(4)=>data_im_in(259),
            data_im_in(5)=>data_im_in(323),
            data_im_in(6)=>data_im_in(387),
            data_im_in(7)=>data_im_in(451),
            data_im_in(8)=>data_im_in(515),
            data_im_in(9)=>data_im_in(579),
            data_im_in(10)=>data_im_in(643),
            data_im_in(11)=>data_im_in(707),
            data_im_in(12)=>data_im_in(771),
            data_im_in(13)=>data_im_in(835),
            data_im_in(14)=>data_im_in(899),
            data_im_in(15)=>data_im_in(963),
            data_im_in(16)=>data_im_in(1027),
            data_im_in(17)=>data_im_in(1091),
            data_im_in(18)=>data_im_in(1155),
            data_im_in(19)=>data_im_in(1219),
            data_im_in(20)=>data_im_in(1283),
            data_im_in(21)=>data_im_in(1347),
            data_im_in(22)=>data_im_in(1411),
            data_im_in(23)=>data_im_in(1475),
            data_im_in(24)=>data_im_in(1539),
            data_im_in(25)=>data_im_in(1603),
            data_im_in(26)=>data_im_in(1667),
            data_im_in(27)=>data_im_in(1731),
            data_im_in(28)=>data_im_in(1795),
            data_im_in(29)=>data_im_in(1859),
            data_im_in(30)=>data_im_in(1923),
            data_im_in(31)=>data_im_in(1987),
            data_re_out=>first_stage_re_out(127 downto 96),
            data_im_out=>first_stage_im_out(127 downto 96)
        );

    ULFFT_PT32_4 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(4),
            data_re_in(1)=>data_re_in(68),
            data_re_in(2)=>data_re_in(132),
            data_re_in(3)=>data_re_in(196),
            data_re_in(4)=>data_re_in(260),
            data_re_in(5)=>data_re_in(324),
            data_re_in(6)=>data_re_in(388),
            data_re_in(7)=>data_re_in(452),
            data_re_in(8)=>data_re_in(516),
            data_re_in(9)=>data_re_in(580),
            data_re_in(10)=>data_re_in(644),
            data_re_in(11)=>data_re_in(708),
            data_re_in(12)=>data_re_in(772),
            data_re_in(13)=>data_re_in(836),
            data_re_in(14)=>data_re_in(900),
            data_re_in(15)=>data_re_in(964),
            data_re_in(16)=>data_re_in(1028),
            data_re_in(17)=>data_re_in(1092),
            data_re_in(18)=>data_re_in(1156),
            data_re_in(19)=>data_re_in(1220),
            data_re_in(20)=>data_re_in(1284),
            data_re_in(21)=>data_re_in(1348),
            data_re_in(22)=>data_re_in(1412),
            data_re_in(23)=>data_re_in(1476),
            data_re_in(24)=>data_re_in(1540),
            data_re_in(25)=>data_re_in(1604),
            data_re_in(26)=>data_re_in(1668),
            data_re_in(27)=>data_re_in(1732),
            data_re_in(28)=>data_re_in(1796),
            data_re_in(29)=>data_re_in(1860),
            data_re_in(30)=>data_re_in(1924),
            data_re_in(31)=>data_re_in(1988),
            data_im_in(0)=>data_im_in(4),
            data_im_in(1)=>data_im_in(68),
            data_im_in(2)=>data_im_in(132),
            data_im_in(3)=>data_im_in(196),
            data_im_in(4)=>data_im_in(260),
            data_im_in(5)=>data_im_in(324),
            data_im_in(6)=>data_im_in(388),
            data_im_in(7)=>data_im_in(452),
            data_im_in(8)=>data_im_in(516),
            data_im_in(9)=>data_im_in(580),
            data_im_in(10)=>data_im_in(644),
            data_im_in(11)=>data_im_in(708),
            data_im_in(12)=>data_im_in(772),
            data_im_in(13)=>data_im_in(836),
            data_im_in(14)=>data_im_in(900),
            data_im_in(15)=>data_im_in(964),
            data_im_in(16)=>data_im_in(1028),
            data_im_in(17)=>data_im_in(1092),
            data_im_in(18)=>data_im_in(1156),
            data_im_in(19)=>data_im_in(1220),
            data_im_in(20)=>data_im_in(1284),
            data_im_in(21)=>data_im_in(1348),
            data_im_in(22)=>data_im_in(1412),
            data_im_in(23)=>data_im_in(1476),
            data_im_in(24)=>data_im_in(1540),
            data_im_in(25)=>data_im_in(1604),
            data_im_in(26)=>data_im_in(1668),
            data_im_in(27)=>data_im_in(1732),
            data_im_in(28)=>data_im_in(1796),
            data_im_in(29)=>data_im_in(1860),
            data_im_in(30)=>data_im_in(1924),
            data_im_in(31)=>data_im_in(1988),
            data_re_out=>first_stage_re_out(159 downto 128),
            data_im_out=>first_stage_im_out(159 downto 128)
        );

    ULFFT_PT32_5 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(5),
            data_re_in(1)=>data_re_in(69),
            data_re_in(2)=>data_re_in(133),
            data_re_in(3)=>data_re_in(197),
            data_re_in(4)=>data_re_in(261),
            data_re_in(5)=>data_re_in(325),
            data_re_in(6)=>data_re_in(389),
            data_re_in(7)=>data_re_in(453),
            data_re_in(8)=>data_re_in(517),
            data_re_in(9)=>data_re_in(581),
            data_re_in(10)=>data_re_in(645),
            data_re_in(11)=>data_re_in(709),
            data_re_in(12)=>data_re_in(773),
            data_re_in(13)=>data_re_in(837),
            data_re_in(14)=>data_re_in(901),
            data_re_in(15)=>data_re_in(965),
            data_re_in(16)=>data_re_in(1029),
            data_re_in(17)=>data_re_in(1093),
            data_re_in(18)=>data_re_in(1157),
            data_re_in(19)=>data_re_in(1221),
            data_re_in(20)=>data_re_in(1285),
            data_re_in(21)=>data_re_in(1349),
            data_re_in(22)=>data_re_in(1413),
            data_re_in(23)=>data_re_in(1477),
            data_re_in(24)=>data_re_in(1541),
            data_re_in(25)=>data_re_in(1605),
            data_re_in(26)=>data_re_in(1669),
            data_re_in(27)=>data_re_in(1733),
            data_re_in(28)=>data_re_in(1797),
            data_re_in(29)=>data_re_in(1861),
            data_re_in(30)=>data_re_in(1925),
            data_re_in(31)=>data_re_in(1989),
            data_im_in(0)=>data_im_in(5),
            data_im_in(1)=>data_im_in(69),
            data_im_in(2)=>data_im_in(133),
            data_im_in(3)=>data_im_in(197),
            data_im_in(4)=>data_im_in(261),
            data_im_in(5)=>data_im_in(325),
            data_im_in(6)=>data_im_in(389),
            data_im_in(7)=>data_im_in(453),
            data_im_in(8)=>data_im_in(517),
            data_im_in(9)=>data_im_in(581),
            data_im_in(10)=>data_im_in(645),
            data_im_in(11)=>data_im_in(709),
            data_im_in(12)=>data_im_in(773),
            data_im_in(13)=>data_im_in(837),
            data_im_in(14)=>data_im_in(901),
            data_im_in(15)=>data_im_in(965),
            data_im_in(16)=>data_im_in(1029),
            data_im_in(17)=>data_im_in(1093),
            data_im_in(18)=>data_im_in(1157),
            data_im_in(19)=>data_im_in(1221),
            data_im_in(20)=>data_im_in(1285),
            data_im_in(21)=>data_im_in(1349),
            data_im_in(22)=>data_im_in(1413),
            data_im_in(23)=>data_im_in(1477),
            data_im_in(24)=>data_im_in(1541),
            data_im_in(25)=>data_im_in(1605),
            data_im_in(26)=>data_im_in(1669),
            data_im_in(27)=>data_im_in(1733),
            data_im_in(28)=>data_im_in(1797),
            data_im_in(29)=>data_im_in(1861),
            data_im_in(30)=>data_im_in(1925),
            data_im_in(31)=>data_im_in(1989),
            data_re_out=>first_stage_re_out(191 downto 160),
            data_im_out=>first_stage_im_out(191 downto 160)
        );

    ULFFT_PT32_6 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(6),
            data_re_in(1)=>data_re_in(70),
            data_re_in(2)=>data_re_in(134),
            data_re_in(3)=>data_re_in(198),
            data_re_in(4)=>data_re_in(262),
            data_re_in(5)=>data_re_in(326),
            data_re_in(6)=>data_re_in(390),
            data_re_in(7)=>data_re_in(454),
            data_re_in(8)=>data_re_in(518),
            data_re_in(9)=>data_re_in(582),
            data_re_in(10)=>data_re_in(646),
            data_re_in(11)=>data_re_in(710),
            data_re_in(12)=>data_re_in(774),
            data_re_in(13)=>data_re_in(838),
            data_re_in(14)=>data_re_in(902),
            data_re_in(15)=>data_re_in(966),
            data_re_in(16)=>data_re_in(1030),
            data_re_in(17)=>data_re_in(1094),
            data_re_in(18)=>data_re_in(1158),
            data_re_in(19)=>data_re_in(1222),
            data_re_in(20)=>data_re_in(1286),
            data_re_in(21)=>data_re_in(1350),
            data_re_in(22)=>data_re_in(1414),
            data_re_in(23)=>data_re_in(1478),
            data_re_in(24)=>data_re_in(1542),
            data_re_in(25)=>data_re_in(1606),
            data_re_in(26)=>data_re_in(1670),
            data_re_in(27)=>data_re_in(1734),
            data_re_in(28)=>data_re_in(1798),
            data_re_in(29)=>data_re_in(1862),
            data_re_in(30)=>data_re_in(1926),
            data_re_in(31)=>data_re_in(1990),
            data_im_in(0)=>data_im_in(6),
            data_im_in(1)=>data_im_in(70),
            data_im_in(2)=>data_im_in(134),
            data_im_in(3)=>data_im_in(198),
            data_im_in(4)=>data_im_in(262),
            data_im_in(5)=>data_im_in(326),
            data_im_in(6)=>data_im_in(390),
            data_im_in(7)=>data_im_in(454),
            data_im_in(8)=>data_im_in(518),
            data_im_in(9)=>data_im_in(582),
            data_im_in(10)=>data_im_in(646),
            data_im_in(11)=>data_im_in(710),
            data_im_in(12)=>data_im_in(774),
            data_im_in(13)=>data_im_in(838),
            data_im_in(14)=>data_im_in(902),
            data_im_in(15)=>data_im_in(966),
            data_im_in(16)=>data_im_in(1030),
            data_im_in(17)=>data_im_in(1094),
            data_im_in(18)=>data_im_in(1158),
            data_im_in(19)=>data_im_in(1222),
            data_im_in(20)=>data_im_in(1286),
            data_im_in(21)=>data_im_in(1350),
            data_im_in(22)=>data_im_in(1414),
            data_im_in(23)=>data_im_in(1478),
            data_im_in(24)=>data_im_in(1542),
            data_im_in(25)=>data_im_in(1606),
            data_im_in(26)=>data_im_in(1670),
            data_im_in(27)=>data_im_in(1734),
            data_im_in(28)=>data_im_in(1798),
            data_im_in(29)=>data_im_in(1862),
            data_im_in(30)=>data_im_in(1926),
            data_im_in(31)=>data_im_in(1990),
            data_re_out=>first_stage_re_out(223 downto 192),
            data_im_out=>first_stage_im_out(223 downto 192)
        );

    ULFFT_PT32_7 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(7),
            data_re_in(1)=>data_re_in(71),
            data_re_in(2)=>data_re_in(135),
            data_re_in(3)=>data_re_in(199),
            data_re_in(4)=>data_re_in(263),
            data_re_in(5)=>data_re_in(327),
            data_re_in(6)=>data_re_in(391),
            data_re_in(7)=>data_re_in(455),
            data_re_in(8)=>data_re_in(519),
            data_re_in(9)=>data_re_in(583),
            data_re_in(10)=>data_re_in(647),
            data_re_in(11)=>data_re_in(711),
            data_re_in(12)=>data_re_in(775),
            data_re_in(13)=>data_re_in(839),
            data_re_in(14)=>data_re_in(903),
            data_re_in(15)=>data_re_in(967),
            data_re_in(16)=>data_re_in(1031),
            data_re_in(17)=>data_re_in(1095),
            data_re_in(18)=>data_re_in(1159),
            data_re_in(19)=>data_re_in(1223),
            data_re_in(20)=>data_re_in(1287),
            data_re_in(21)=>data_re_in(1351),
            data_re_in(22)=>data_re_in(1415),
            data_re_in(23)=>data_re_in(1479),
            data_re_in(24)=>data_re_in(1543),
            data_re_in(25)=>data_re_in(1607),
            data_re_in(26)=>data_re_in(1671),
            data_re_in(27)=>data_re_in(1735),
            data_re_in(28)=>data_re_in(1799),
            data_re_in(29)=>data_re_in(1863),
            data_re_in(30)=>data_re_in(1927),
            data_re_in(31)=>data_re_in(1991),
            data_im_in(0)=>data_im_in(7),
            data_im_in(1)=>data_im_in(71),
            data_im_in(2)=>data_im_in(135),
            data_im_in(3)=>data_im_in(199),
            data_im_in(4)=>data_im_in(263),
            data_im_in(5)=>data_im_in(327),
            data_im_in(6)=>data_im_in(391),
            data_im_in(7)=>data_im_in(455),
            data_im_in(8)=>data_im_in(519),
            data_im_in(9)=>data_im_in(583),
            data_im_in(10)=>data_im_in(647),
            data_im_in(11)=>data_im_in(711),
            data_im_in(12)=>data_im_in(775),
            data_im_in(13)=>data_im_in(839),
            data_im_in(14)=>data_im_in(903),
            data_im_in(15)=>data_im_in(967),
            data_im_in(16)=>data_im_in(1031),
            data_im_in(17)=>data_im_in(1095),
            data_im_in(18)=>data_im_in(1159),
            data_im_in(19)=>data_im_in(1223),
            data_im_in(20)=>data_im_in(1287),
            data_im_in(21)=>data_im_in(1351),
            data_im_in(22)=>data_im_in(1415),
            data_im_in(23)=>data_im_in(1479),
            data_im_in(24)=>data_im_in(1543),
            data_im_in(25)=>data_im_in(1607),
            data_im_in(26)=>data_im_in(1671),
            data_im_in(27)=>data_im_in(1735),
            data_im_in(28)=>data_im_in(1799),
            data_im_in(29)=>data_im_in(1863),
            data_im_in(30)=>data_im_in(1927),
            data_im_in(31)=>data_im_in(1991),
            data_re_out=>first_stage_re_out(255 downto 224),
            data_im_out=>first_stage_im_out(255 downto 224)
        );

    ULFFT_PT32_8 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(8),
            data_re_in(1)=>data_re_in(72),
            data_re_in(2)=>data_re_in(136),
            data_re_in(3)=>data_re_in(200),
            data_re_in(4)=>data_re_in(264),
            data_re_in(5)=>data_re_in(328),
            data_re_in(6)=>data_re_in(392),
            data_re_in(7)=>data_re_in(456),
            data_re_in(8)=>data_re_in(520),
            data_re_in(9)=>data_re_in(584),
            data_re_in(10)=>data_re_in(648),
            data_re_in(11)=>data_re_in(712),
            data_re_in(12)=>data_re_in(776),
            data_re_in(13)=>data_re_in(840),
            data_re_in(14)=>data_re_in(904),
            data_re_in(15)=>data_re_in(968),
            data_re_in(16)=>data_re_in(1032),
            data_re_in(17)=>data_re_in(1096),
            data_re_in(18)=>data_re_in(1160),
            data_re_in(19)=>data_re_in(1224),
            data_re_in(20)=>data_re_in(1288),
            data_re_in(21)=>data_re_in(1352),
            data_re_in(22)=>data_re_in(1416),
            data_re_in(23)=>data_re_in(1480),
            data_re_in(24)=>data_re_in(1544),
            data_re_in(25)=>data_re_in(1608),
            data_re_in(26)=>data_re_in(1672),
            data_re_in(27)=>data_re_in(1736),
            data_re_in(28)=>data_re_in(1800),
            data_re_in(29)=>data_re_in(1864),
            data_re_in(30)=>data_re_in(1928),
            data_re_in(31)=>data_re_in(1992),
            data_im_in(0)=>data_im_in(8),
            data_im_in(1)=>data_im_in(72),
            data_im_in(2)=>data_im_in(136),
            data_im_in(3)=>data_im_in(200),
            data_im_in(4)=>data_im_in(264),
            data_im_in(5)=>data_im_in(328),
            data_im_in(6)=>data_im_in(392),
            data_im_in(7)=>data_im_in(456),
            data_im_in(8)=>data_im_in(520),
            data_im_in(9)=>data_im_in(584),
            data_im_in(10)=>data_im_in(648),
            data_im_in(11)=>data_im_in(712),
            data_im_in(12)=>data_im_in(776),
            data_im_in(13)=>data_im_in(840),
            data_im_in(14)=>data_im_in(904),
            data_im_in(15)=>data_im_in(968),
            data_im_in(16)=>data_im_in(1032),
            data_im_in(17)=>data_im_in(1096),
            data_im_in(18)=>data_im_in(1160),
            data_im_in(19)=>data_im_in(1224),
            data_im_in(20)=>data_im_in(1288),
            data_im_in(21)=>data_im_in(1352),
            data_im_in(22)=>data_im_in(1416),
            data_im_in(23)=>data_im_in(1480),
            data_im_in(24)=>data_im_in(1544),
            data_im_in(25)=>data_im_in(1608),
            data_im_in(26)=>data_im_in(1672),
            data_im_in(27)=>data_im_in(1736),
            data_im_in(28)=>data_im_in(1800),
            data_im_in(29)=>data_im_in(1864),
            data_im_in(30)=>data_im_in(1928),
            data_im_in(31)=>data_im_in(1992),
            data_re_out=>first_stage_re_out(287 downto 256),
            data_im_out=>first_stage_im_out(287 downto 256)
        );

    ULFFT_PT32_9 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(9),
            data_re_in(1)=>data_re_in(73),
            data_re_in(2)=>data_re_in(137),
            data_re_in(3)=>data_re_in(201),
            data_re_in(4)=>data_re_in(265),
            data_re_in(5)=>data_re_in(329),
            data_re_in(6)=>data_re_in(393),
            data_re_in(7)=>data_re_in(457),
            data_re_in(8)=>data_re_in(521),
            data_re_in(9)=>data_re_in(585),
            data_re_in(10)=>data_re_in(649),
            data_re_in(11)=>data_re_in(713),
            data_re_in(12)=>data_re_in(777),
            data_re_in(13)=>data_re_in(841),
            data_re_in(14)=>data_re_in(905),
            data_re_in(15)=>data_re_in(969),
            data_re_in(16)=>data_re_in(1033),
            data_re_in(17)=>data_re_in(1097),
            data_re_in(18)=>data_re_in(1161),
            data_re_in(19)=>data_re_in(1225),
            data_re_in(20)=>data_re_in(1289),
            data_re_in(21)=>data_re_in(1353),
            data_re_in(22)=>data_re_in(1417),
            data_re_in(23)=>data_re_in(1481),
            data_re_in(24)=>data_re_in(1545),
            data_re_in(25)=>data_re_in(1609),
            data_re_in(26)=>data_re_in(1673),
            data_re_in(27)=>data_re_in(1737),
            data_re_in(28)=>data_re_in(1801),
            data_re_in(29)=>data_re_in(1865),
            data_re_in(30)=>data_re_in(1929),
            data_re_in(31)=>data_re_in(1993),
            data_im_in(0)=>data_im_in(9),
            data_im_in(1)=>data_im_in(73),
            data_im_in(2)=>data_im_in(137),
            data_im_in(3)=>data_im_in(201),
            data_im_in(4)=>data_im_in(265),
            data_im_in(5)=>data_im_in(329),
            data_im_in(6)=>data_im_in(393),
            data_im_in(7)=>data_im_in(457),
            data_im_in(8)=>data_im_in(521),
            data_im_in(9)=>data_im_in(585),
            data_im_in(10)=>data_im_in(649),
            data_im_in(11)=>data_im_in(713),
            data_im_in(12)=>data_im_in(777),
            data_im_in(13)=>data_im_in(841),
            data_im_in(14)=>data_im_in(905),
            data_im_in(15)=>data_im_in(969),
            data_im_in(16)=>data_im_in(1033),
            data_im_in(17)=>data_im_in(1097),
            data_im_in(18)=>data_im_in(1161),
            data_im_in(19)=>data_im_in(1225),
            data_im_in(20)=>data_im_in(1289),
            data_im_in(21)=>data_im_in(1353),
            data_im_in(22)=>data_im_in(1417),
            data_im_in(23)=>data_im_in(1481),
            data_im_in(24)=>data_im_in(1545),
            data_im_in(25)=>data_im_in(1609),
            data_im_in(26)=>data_im_in(1673),
            data_im_in(27)=>data_im_in(1737),
            data_im_in(28)=>data_im_in(1801),
            data_im_in(29)=>data_im_in(1865),
            data_im_in(30)=>data_im_in(1929),
            data_im_in(31)=>data_im_in(1993),
            data_re_out=>first_stage_re_out(319 downto 288),
            data_im_out=>first_stage_im_out(319 downto 288)
        );

    ULFFT_PT32_10 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(10),
            data_re_in(1)=>data_re_in(74),
            data_re_in(2)=>data_re_in(138),
            data_re_in(3)=>data_re_in(202),
            data_re_in(4)=>data_re_in(266),
            data_re_in(5)=>data_re_in(330),
            data_re_in(6)=>data_re_in(394),
            data_re_in(7)=>data_re_in(458),
            data_re_in(8)=>data_re_in(522),
            data_re_in(9)=>data_re_in(586),
            data_re_in(10)=>data_re_in(650),
            data_re_in(11)=>data_re_in(714),
            data_re_in(12)=>data_re_in(778),
            data_re_in(13)=>data_re_in(842),
            data_re_in(14)=>data_re_in(906),
            data_re_in(15)=>data_re_in(970),
            data_re_in(16)=>data_re_in(1034),
            data_re_in(17)=>data_re_in(1098),
            data_re_in(18)=>data_re_in(1162),
            data_re_in(19)=>data_re_in(1226),
            data_re_in(20)=>data_re_in(1290),
            data_re_in(21)=>data_re_in(1354),
            data_re_in(22)=>data_re_in(1418),
            data_re_in(23)=>data_re_in(1482),
            data_re_in(24)=>data_re_in(1546),
            data_re_in(25)=>data_re_in(1610),
            data_re_in(26)=>data_re_in(1674),
            data_re_in(27)=>data_re_in(1738),
            data_re_in(28)=>data_re_in(1802),
            data_re_in(29)=>data_re_in(1866),
            data_re_in(30)=>data_re_in(1930),
            data_re_in(31)=>data_re_in(1994),
            data_im_in(0)=>data_im_in(10),
            data_im_in(1)=>data_im_in(74),
            data_im_in(2)=>data_im_in(138),
            data_im_in(3)=>data_im_in(202),
            data_im_in(4)=>data_im_in(266),
            data_im_in(5)=>data_im_in(330),
            data_im_in(6)=>data_im_in(394),
            data_im_in(7)=>data_im_in(458),
            data_im_in(8)=>data_im_in(522),
            data_im_in(9)=>data_im_in(586),
            data_im_in(10)=>data_im_in(650),
            data_im_in(11)=>data_im_in(714),
            data_im_in(12)=>data_im_in(778),
            data_im_in(13)=>data_im_in(842),
            data_im_in(14)=>data_im_in(906),
            data_im_in(15)=>data_im_in(970),
            data_im_in(16)=>data_im_in(1034),
            data_im_in(17)=>data_im_in(1098),
            data_im_in(18)=>data_im_in(1162),
            data_im_in(19)=>data_im_in(1226),
            data_im_in(20)=>data_im_in(1290),
            data_im_in(21)=>data_im_in(1354),
            data_im_in(22)=>data_im_in(1418),
            data_im_in(23)=>data_im_in(1482),
            data_im_in(24)=>data_im_in(1546),
            data_im_in(25)=>data_im_in(1610),
            data_im_in(26)=>data_im_in(1674),
            data_im_in(27)=>data_im_in(1738),
            data_im_in(28)=>data_im_in(1802),
            data_im_in(29)=>data_im_in(1866),
            data_im_in(30)=>data_im_in(1930),
            data_im_in(31)=>data_im_in(1994),
            data_re_out=>first_stage_re_out(351 downto 320),
            data_im_out=>first_stage_im_out(351 downto 320)
        );

    ULFFT_PT32_11 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(11),
            data_re_in(1)=>data_re_in(75),
            data_re_in(2)=>data_re_in(139),
            data_re_in(3)=>data_re_in(203),
            data_re_in(4)=>data_re_in(267),
            data_re_in(5)=>data_re_in(331),
            data_re_in(6)=>data_re_in(395),
            data_re_in(7)=>data_re_in(459),
            data_re_in(8)=>data_re_in(523),
            data_re_in(9)=>data_re_in(587),
            data_re_in(10)=>data_re_in(651),
            data_re_in(11)=>data_re_in(715),
            data_re_in(12)=>data_re_in(779),
            data_re_in(13)=>data_re_in(843),
            data_re_in(14)=>data_re_in(907),
            data_re_in(15)=>data_re_in(971),
            data_re_in(16)=>data_re_in(1035),
            data_re_in(17)=>data_re_in(1099),
            data_re_in(18)=>data_re_in(1163),
            data_re_in(19)=>data_re_in(1227),
            data_re_in(20)=>data_re_in(1291),
            data_re_in(21)=>data_re_in(1355),
            data_re_in(22)=>data_re_in(1419),
            data_re_in(23)=>data_re_in(1483),
            data_re_in(24)=>data_re_in(1547),
            data_re_in(25)=>data_re_in(1611),
            data_re_in(26)=>data_re_in(1675),
            data_re_in(27)=>data_re_in(1739),
            data_re_in(28)=>data_re_in(1803),
            data_re_in(29)=>data_re_in(1867),
            data_re_in(30)=>data_re_in(1931),
            data_re_in(31)=>data_re_in(1995),
            data_im_in(0)=>data_im_in(11),
            data_im_in(1)=>data_im_in(75),
            data_im_in(2)=>data_im_in(139),
            data_im_in(3)=>data_im_in(203),
            data_im_in(4)=>data_im_in(267),
            data_im_in(5)=>data_im_in(331),
            data_im_in(6)=>data_im_in(395),
            data_im_in(7)=>data_im_in(459),
            data_im_in(8)=>data_im_in(523),
            data_im_in(9)=>data_im_in(587),
            data_im_in(10)=>data_im_in(651),
            data_im_in(11)=>data_im_in(715),
            data_im_in(12)=>data_im_in(779),
            data_im_in(13)=>data_im_in(843),
            data_im_in(14)=>data_im_in(907),
            data_im_in(15)=>data_im_in(971),
            data_im_in(16)=>data_im_in(1035),
            data_im_in(17)=>data_im_in(1099),
            data_im_in(18)=>data_im_in(1163),
            data_im_in(19)=>data_im_in(1227),
            data_im_in(20)=>data_im_in(1291),
            data_im_in(21)=>data_im_in(1355),
            data_im_in(22)=>data_im_in(1419),
            data_im_in(23)=>data_im_in(1483),
            data_im_in(24)=>data_im_in(1547),
            data_im_in(25)=>data_im_in(1611),
            data_im_in(26)=>data_im_in(1675),
            data_im_in(27)=>data_im_in(1739),
            data_im_in(28)=>data_im_in(1803),
            data_im_in(29)=>data_im_in(1867),
            data_im_in(30)=>data_im_in(1931),
            data_im_in(31)=>data_im_in(1995),
            data_re_out=>first_stage_re_out(383 downto 352),
            data_im_out=>first_stage_im_out(383 downto 352)
        );

    ULFFT_PT32_12 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(12),
            data_re_in(1)=>data_re_in(76),
            data_re_in(2)=>data_re_in(140),
            data_re_in(3)=>data_re_in(204),
            data_re_in(4)=>data_re_in(268),
            data_re_in(5)=>data_re_in(332),
            data_re_in(6)=>data_re_in(396),
            data_re_in(7)=>data_re_in(460),
            data_re_in(8)=>data_re_in(524),
            data_re_in(9)=>data_re_in(588),
            data_re_in(10)=>data_re_in(652),
            data_re_in(11)=>data_re_in(716),
            data_re_in(12)=>data_re_in(780),
            data_re_in(13)=>data_re_in(844),
            data_re_in(14)=>data_re_in(908),
            data_re_in(15)=>data_re_in(972),
            data_re_in(16)=>data_re_in(1036),
            data_re_in(17)=>data_re_in(1100),
            data_re_in(18)=>data_re_in(1164),
            data_re_in(19)=>data_re_in(1228),
            data_re_in(20)=>data_re_in(1292),
            data_re_in(21)=>data_re_in(1356),
            data_re_in(22)=>data_re_in(1420),
            data_re_in(23)=>data_re_in(1484),
            data_re_in(24)=>data_re_in(1548),
            data_re_in(25)=>data_re_in(1612),
            data_re_in(26)=>data_re_in(1676),
            data_re_in(27)=>data_re_in(1740),
            data_re_in(28)=>data_re_in(1804),
            data_re_in(29)=>data_re_in(1868),
            data_re_in(30)=>data_re_in(1932),
            data_re_in(31)=>data_re_in(1996),
            data_im_in(0)=>data_im_in(12),
            data_im_in(1)=>data_im_in(76),
            data_im_in(2)=>data_im_in(140),
            data_im_in(3)=>data_im_in(204),
            data_im_in(4)=>data_im_in(268),
            data_im_in(5)=>data_im_in(332),
            data_im_in(6)=>data_im_in(396),
            data_im_in(7)=>data_im_in(460),
            data_im_in(8)=>data_im_in(524),
            data_im_in(9)=>data_im_in(588),
            data_im_in(10)=>data_im_in(652),
            data_im_in(11)=>data_im_in(716),
            data_im_in(12)=>data_im_in(780),
            data_im_in(13)=>data_im_in(844),
            data_im_in(14)=>data_im_in(908),
            data_im_in(15)=>data_im_in(972),
            data_im_in(16)=>data_im_in(1036),
            data_im_in(17)=>data_im_in(1100),
            data_im_in(18)=>data_im_in(1164),
            data_im_in(19)=>data_im_in(1228),
            data_im_in(20)=>data_im_in(1292),
            data_im_in(21)=>data_im_in(1356),
            data_im_in(22)=>data_im_in(1420),
            data_im_in(23)=>data_im_in(1484),
            data_im_in(24)=>data_im_in(1548),
            data_im_in(25)=>data_im_in(1612),
            data_im_in(26)=>data_im_in(1676),
            data_im_in(27)=>data_im_in(1740),
            data_im_in(28)=>data_im_in(1804),
            data_im_in(29)=>data_im_in(1868),
            data_im_in(30)=>data_im_in(1932),
            data_im_in(31)=>data_im_in(1996),
            data_re_out=>first_stage_re_out(415 downto 384),
            data_im_out=>first_stage_im_out(415 downto 384)
        );

    ULFFT_PT32_13 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(13),
            data_re_in(1)=>data_re_in(77),
            data_re_in(2)=>data_re_in(141),
            data_re_in(3)=>data_re_in(205),
            data_re_in(4)=>data_re_in(269),
            data_re_in(5)=>data_re_in(333),
            data_re_in(6)=>data_re_in(397),
            data_re_in(7)=>data_re_in(461),
            data_re_in(8)=>data_re_in(525),
            data_re_in(9)=>data_re_in(589),
            data_re_in(10)=>data_re_in(653),
            data_re_in(11)=>data_re_in(717),
            data_re_in(12)=>data_re_in(781),
            data_re_in(13)=>data_re_in(845),
            data_re_in(14)=>data_re_in(909),
            data_re_in(15)=>data_re_in(973),
            data_re_in(16)=>data_re_in(1037),
            data_re_in(17)=>data_re_in(1101),
            data_re_in(18)=>data_re_in(1165),
            data_re_in(19)=>data_re_in(1229),
            data_re_in(20)=>data_re_in(1293),
            data_re_in(21)=>data_re_in(1357),
            data_re_in(22)=>data_re_in(1421),
            data_re_in(23)=>data_re_in(1485),
            data_re_in(24)=>data_re_in(1549),
            data_re_in(25)=>data_re_in(1613),
            data_re_in(26)=>data_re_in(1677),
            data_re_in(27)=>data_re_in(1741),
            data_re_in(28)=>data_re_in(1805),
            data_re_in(29)=>data_re_in(1869),
            data_re_in(30)=>data_re_in(1933),
            data_re_in(31)=>data_re_in(1997),
            data_im_in(0)=>data_im_in(13),
            data_im_in(1)=>data_im_in(77),
            data_im_in(2)=>data_im_in(141),
            data_im_in(3)=>data_im_in(205),
            data_im_in(4)=>data_im_in(269),
            data_im_in(5)=>data_im_in(333),
            data_im_in(6)=>data_im_in(397),
            data_im_in(7)=>data_im_in(461),
            data_im_in(8)=>data_im_in(525),
            data_im_in(9)=>data_im_in(589),
            data_im_in(10)=>data_im_in(653),
            data_im_in(11)=>data_im_in(717),
            data_im_in(12)=>data_im_in(781),
            data_im_in(13)=>data_im_in(845),
            data_im_in(14)=>data_im_in(909),
            data_im_in(15)=>data_im_in(973),
            data_im_in(16)=>data_im_in(1037),
            data_im_in(17)=>data_im_in(1101),
            data_im_in(18)=>data_im_in(1165),
            data_im_in(19)=>data_im_in(1229),
            data_im_in(20)=>data_im_in(1293),
            data_im_in(21)=>data_im_in(1357),
            data_im_in(22)=>data_im_in(1421),
            data_im_in(23)=>data_im_in(1485),
            data_im_in(24)=>data_im_in(1549),
            data_im_in(25)=>data_im_in(1613),
            data_im_in(26)=>data_im_in(1677),
            data_im_in(27)=>data_im_in(1741),
            data_im_in(28)=>data_im_in(1805),
            data_im_in(29)=>data_im_in(1869),
            data_im_in(30)=>data_im_in(1933),
            data_im_in(31)=>data_im_in(1997),
            data_re_out=>first_stage_re_out(447 downto 416),
            data_im_out=>first_stage_im_out(447 downto 416)
        );

    ULFFT_PT32_14 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(14),
            data_re_in(1)=>data_re_in(78),
            data_re_in(2)=>data_re_in(142),
            data_re_in(3)=>data_re_in(206),
            data_re_in(4)=>data_re_in(270),
            data_re_in(5)=>data_re_in(334),
            data_re_in(6)=>data_re_in(398),
            data_re_in(7)=>data_re_in(462),
            data_re_in(8)=>data_re_in(526),
            data_re_in(9)=>data_re_in(590),
            data_re_in(10)=>data_re_in(654),
            data_re_in(11)=>data_re_in(718),
            data_re_in(12)=>data_re_in(782),
            data_re_in(13)=>data_re_in(846),
            data_re_in(14)=>data_re_in(910),
            data_re_in(15)=>data_re_in(974),
            data_re_in(16)=>data_re_in(1038),
            data_re_in(17)=>data_re_in(1102),
            data_re_in(18)=>data_re_in(1166),
            data_re_in(19)=>data_re_in(1230),
            data_re_in(20)=>data_re_in(1294),
            data_re_in(21)=>data_re_in(1358),
            data_re_in(22)=>data_re_in(1422),
            data_re_in(23)=>data_re_in(1486),
            data_re_in(24)=>data_re_in(1550),
            data_re_in(25)=>data_re_in(1614),
            data_re_in(26)=>data_re_in(1678),
            data_re_in(27)=>data_re_in(1742),
            data_re_in(28)=>data_re_in(1806),
            data_re_in(29)=>data_re_in(1870),
            data_re_in(30)=>data_re_in(1934),
            data_re_in(31)=>data_re_in(1998),
            data_im_in(0)=>data_im_in(14),
            data_im_in(1)=>data_im_in(78),
            data_im_in(2)=>data_im_in(142),
            data_im_in(3)=>data_im_in(206),
            data_im_in(4)=>data_im_in(270),
            data_im_in(5)=>data_im_in(334),
            data_im_in(6)=>data_im_in(398),
            data_im_in(7)=>data_im_in(462),
            data_im_in(8)=>data_im_in(526),
            data_im_in(9)=>data_im_in(590),
            data_im_in(10)=>data_im_in(654),
            data_im_in(11)=>data_im_in(718),
            data_im_in(12)=>data_im_in(782),
            data_im_in(13)=>data_im_in(846),
            data_im_in(14)=>data_im_in(910),
            data_im_in(15)=>data_im_in(974),
            data_im_in(16)=>data_im_in(1038),
            data_im_in(17)=>data_im_in(1102),
            data_im_in(18)=>data_im_in(1166),
            data_im_in(19)=>data_im_in(1230),
            data_im_in(20)=>data_im_in(1294),
            data_im_in(21)=>data_im_in(1358),
            data_im_in(22)=>data_im_in(1422),
            data_im_in(23)=>data_im_in(1486),
            data_im_in(24)=>data_im_in(1550),
            data_im_in(25)=>data_im_in(1614),
            data_im_in(26)=>data_im_in(1678),
            data_im_in(27)=>data_im_in(1742),
            data_im_in(28)=>data_im_in(1806),
            data_im_in(29)=>data_im_in(1870),
            data_im_in(30)=>data_im_in(1934),
            data_im_in(31)=>data_im_in(1998),
            data_re_out=>first_stage_re_out(479 downto 448),
            data_im_out=>first_stage_im_out(479 downto 448)
        );

    ULFFT_PT32_15 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(15),
            data_re_in(1)=>data_re_in(79),
            data_re_in(2)=>data_re_in(143),
            data_re_in(3)=>data_re_in(207),
            data_re_in(4)=>data_re_in(271),
            data_re_in(5)=>data_re_in(335),
            data_re_in(6)=>data_re_in(399),
            data_re_in(7)=>data_re_in(463),
            data_re_in(8)=>data_re_in(527),
            data_re_in(9)=>data_re_in(591),
            data_re_in(10)=>data_re_in(655),
            data_re_in(11)=>data_re_in(719),
            data_re_in(12)=>data_re_in(783),
            data_re_in(13)=>data_re_in(847),
            data_re_in(14)=>data_re_in(911),
            data_re_in(15)=>data_re_in(975),
            data_re_in(16)=>data_re_in(1039),
            data_re_in(17)=>data_re_in(1103),
            data_re_in(18)=>data_re_in(1167),
            data_re_in(19)=>data_re_in(1231),
            data_re_in(20)=>data_re_in(1295),
            data_re_in(21)=>data_re_in(1359),
            data_re_in(22)=>data_re_in(1423),
            data_re_in(23)=>data_re_in(1487),
            data_re_in(24)=>data_re_in(1551),
            data_re_in(25)=>data_re_in(1615),
            data_re_in(26)=>data_re_in(1679),
            data_re_in(27)=>data_re_in(1743),
            data_re_in(28)=>data_re_in(1807),
            data_re_in(29)=>data_re_in(1871),
            data_re_in(30)=>data_re_in(1935),
            data_re_in(31)=>data_re_in(1999),
            data_im_in(0)=>data_im_in(15),
            data_im_in(1)=>data_im_in(79),
            data_im_in(2)=>data_im_in(143),
            data_im_in(3)=>data_im_in(207),
            data_im_in(4)=>data_im_in(271),
            data_im_in(5)=>data_im_in(335),
            data_im_in(6)=>data_im_in(399),
            data_im_in(7)=>data_im_in(463),
            data_im_in(8)=>data_im_in(527),
            data_im_in(9)=>data_im_in(591),
            data_im_in(10)=>data_im_in(655),
            data_im_in(11)=>data_im_in(719),
            data_im_in(12)=>data_im_in(783),
            data_im_in(13)=>data_im_in(847),
            data_im_in(14)=>data_im_in(911),
            data_im_in(15)=>data_im_in(975),
            data_im_in(16)=>data_im_in(1039),
            data_im_in(17)=>data_im_in(1103),
            data_im_in(18)=>data_im_in(1167),
            data_im_in(19)=>data_im_in(1231),
            data_im_in(20)=>data_im_in(1295),
            data_im_in(21)=>data_im_in(1359),
            data_im_in(22)=>data_im_in(1423),
            data_im_in(23)=>data_im_in(1487),
            data_im_in(24)=>data_im_in(1551),
            data_im_in(25)=>data_im_in(1615),
            data_im_in(26)=>data_im_in(1679),
            data_im_in(27)=>data_im_in(1743),
            data_im_in(28)=>data_im_in(1807),
            data_im_in(29)=>data_im_in(1871),
            data_im_in(30)=>data_im_in(1935),
            data_im_in(31)=>data_im_in(1999),
            data_re_out=>first_stage_re_out(511 downto 480),
            data_im_out=>first_stage_im_out(511 downto 480)
        );

    ULFFT_PT32_16 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(16),
            data_re_in(1)=>data_re_in(80),
            data_re_in(2)=>data_re_in(144),
            data_re_in(3)=>data_re_in(208),
            data_re_in(4)=>data_re_in(272),
            data_re_in(5)=>data_re_in(336),
            data_re_in(6)=>data_re_in(400),
            data_re_in(7)=>data_re_in(464),
            data_re_in(8)=>data_re_in(528),
            data_re_in(9)=>data_re_in(592),
            data_re_in(10)=>data_re_in(656),
            data_re_in(11)=>data_re_in(720),
            data_re_in(12)=>data_re_in(784),
            data_re_in(13)=>data_re_in(848),
            data_re_in(14)=>data_re_in(912),
            data_re_in(15)=>data_re_in(976),
            data_re_in(16)=>data_re_in(1040),
            data_re_in(17)=>data_re_in(1104),
            data_re_in(18)=>data_re_in(1168),
            data_re_in(19)=>data_re_in(1232),
            data_re_in(20)=>data_re_in(1296),
            data_re_in(21)=>data_re_in(1360),
            data_re_in(22)=>data_re_in(1424),
            data_re_in(23)=>data_re_in(1488),
            data_re_in(24)=>data_re_in(1552),
            data_re_in(25)=>data_re_in(1616),
            data_re_in(26)=>data_re_in(1680),
            data_re_in(27)=>data_re_in(1744),
            data_re_in(28)=>data_re_in(1808),
            data_re_in(29)=>data_re_in(1872),
            data_re_in(30)=>data_re_in(1936),
            data_re_in(31)=>data_re_in(2000),
            data_im_in(0)=>data_im_in(16),
            data_im_in(1)=>data_im_in(80),
            data_im_in(2)=>data_im_in(144),
            data_im_in(3)=>data_im_in(208),
            data_im_in(4)=>data_im_in(272),
            data_im_in(5)=>data_im_in(336),
            data_im_in(6)=>data_im_in(400),
            data_im_in(7)=>data_im_in(464),
            data_im_in(8)=>data_im_in(528),
            data_im_in(9)=>data_im_in(592),
            data_im_in(10)=>data_im_in(656),
            data_im_in(11)=>data_im_in(720),
            data_im_in(12)=>data_im_in(784),
            data_im_in(13)=>data_im_in(848),
            data_im_in(14)=>data_im_in(912),
            data_im_in(15)=>data_im_in(976),
            data_im_in(16)=>data_im_in(1040),
            data_im_in(17)=>data_im_in(1104),
            data_im_in(18)=>data_im_in(1168),
            data_im_in(19)=>data_im_in(1232),
            data_im_in(20)=>data_im_in(1296),
            data_im_in(21)=>data_im_in(1360),
            data_im_in(22)=>data_im_in(1424),
            data_im_in(23)=>data_im_in(1488),
            data_im_in(24)=>data_im_in(1552),
            data_im_in(25)=>data_im_in(1616),
            data_im_in(26)=>data_im_in(1680),
            data_im_in(27)=>data_im_in(1744),
            data_im_in(28)=>data_im_in(1808),
            data_im_in(29)=>data_im_in(1872),
            data_im_in(30)=>data_im_in(1936),
            data_im_in(31)=>data_im_in(2000),
            data_re_out=>first_stage_re_out(543 downto 512),
            data_im_out=>first_stage_im_out(543 downto 512)
        );

    ULFFT_PT32_17 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(17),
            data_re_in(1)=>data_re_in(81),
            data_re_in(2)=>data_re_in(145),
            data_re_in(3)=>data_re_in(209),
            data_re_in(4)=>data_re_in(273),
            data_re_in(5)=>data_re_in(337),
            data_re_in(6)=>data_re_in(401),
            data_re_in(7)=>data_re_in(465),
            data_re_in(8)=>data_re_in(529),
            data_re_in(9)=>data_re_in(593),
            data_re_in(10)=>data_re_in(657),
            data_re_in(11)=>data_re_in(721),
            data_re_in(12)=>data_re_in(785),
            data_re_in(13)=>data_re_in(849),
            data_re_in(14)=>data_re_in(913),
            data_re_in(15)=>data_re_in(977),
            data_re_in(16)=>data_re_in(1041),
            data_re_in(17)=>data_re_in(1105),
            data_re_in(18)=>data_re_in(1169),
            data_re_in(19)=>data_re_in(1233),
            data_re_in(20)=>data_re_in(1297),
            data_re_in(21)=>data_re_in(1361),
            data_re_in(22)=>data_re_in(1425),
            data_re_in(23)=>data_re_in(1489),
            data_re_in(24)=>data_re_in(1553),
            data_re_in(25)=>data_re_in(1617),
            data_re_in(26)=>data_re_in(1681),
            data_re_in(27)=>data_re_in(1745),
            data_re_in(28)=>data_re_in(1809),
            data_re_in(29)=>data_re_in(1873),
            data_re_in(30)=>data_re_in(1937),
            data_re_in(31)=>data_re_in(2001),
            data_im_in(0)=>data_im_in(17),
            data_im_in(1)=>data_im_in(81),
            data_im_in(2)=>data_im_in(145),
            data_im_in(3)=>data_im_in(209),
            data_im_in(4)=>data_im_in(273),
            data_im_in(5)=>data_im_in(337),
            data_im_in(6)=>data_im_in(401),
            data_im_in(7)=>data_im_in(465),
            data_im_in(8)=>data_im_in(529),
            data_im_in(9)=>data_im_in(593),
            data_im_in(10)=>data_im_in(657),
            data_im_in(11)=>data_im_in(721),
            data_im_in(12)=>data_im_in(785),
            data_im_in(13)=>data_im_in(849),
            data_im_in(14)=>data_im_in(913),
            data_im_in(15)=>data_im_in(977),
            data_im_in(16)=>data_im_in(1041),
            data_im_in(17)=>data_im_in(1105),
            data_im_in(18)=>data_im_in(1169),
            data_im_in(19)=>data_im_in(1233),
            data_im_in(20)=>data_im_in(1297),
            data_im_in(21)=>data_im_in(1361),
            data_im_in(22)=>data_im_in(1425),
            data_im_in(23)=>data_im_in(1489),
            data_im_in(24)=>data_im_in(1553),
            data_im_in(25)=>data_im_in(1617),
            data_im_in(26)=>data_im_in(1681),
            data_im_in(27)=>data_im_in(1745),
            data_im_in(28)=>data_im_in(1809),
            data_im_in(29)=>data_im_in(1873),
            data_im_in(30)=>data_im_in(1937),
            data_im_in(31)=>data_im_in(2001),
            data_re_out=>first_stage_re_out(575 downto 544),
            data_im_out=>first_stage_im_out(575 downto 544)
        );

    ULFFT_PT32_18 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(18),
            data_re_in(1)=>data_re_in(82),
            data_re_in(2)=>data_re_in(146),
            data_re_in(3)=>data_re_in(210),
            data_re_in(4)=>data_re_in(274),
            data_re_in(5)=>data_re_in(338),
            data_re_in(6)=>data_re_in(402),
            data_re_in(7)=>data_re_in(466),
            data_re_in(8)=>data_re_in(530),
            data_re_in(9)=>data_re_in(594),
            data_re_in(10)=>data_re_in(658),
            data_re_in(11)=>data_re_in(722),
            data_re_in(12)=>data_re_in(786),
            data_re_in(13)=>data_re_in(850),
            data_re_in(14)=>data_re_in(914),
            data_re_in(15)=>data_re_in(978),
            data_re_in(16)=>data_re_in(1042),
            data_re_in(17)=>data_re_in(1106),
            data_re_in(18)=>data_re_in(1170),
            data_re_in(19)=>data_re_in(1234),
            data_re_in(20)=>data_re_in(1298),
            data_re_in(21)=>data_re_in(1362),
            data_re_in(22)=>data_re_in(1426),
            data_re_in(23)=>data_re_in(1490),
            data_re_in(24)=>data_re_in(1554),
            data_re_in(25)=>data_re_in(1618),
            data_re_in(26)=>data_re_in(1682),
            data_re_in(27)=>data_re_in(1746),
            data_re_in(28)=>data_re_in(1810),
            data_re_in(29)=>data_re_in(1874),
            data_re_in(30)=>data_re_in(1938),
            data_re_in(31)=>data_re_in(2002),
            data_im_in(0)=>data_im_in(18),
            data_im_in(1)=>data_im_in(82),
            data_im_in(2)=>data_im_in(146),
            data_im_in(3)=>data_im_in(210),
            data_im_in(4)=>data_im_in(274),
            data_im_in(5)=>data_im_in(338),
            data_im_in(6)=>data_im_in(402),
            data_im_in(7)=>data_im_in(466),
            data_im_in(8)=>data_im_in(530),
            data_im_in(9)=>data_im_in(594),
            data_im_in(10)=>data_im_in(658),
            data_im_in(11)=>data_im_in(722),
            data_im_in(12)=>data_im_in(786),
            data_im_in(13)=>data_im_in(850),
            data_im_in(14)=>data_im_in(914),
            data_im_in(15)=>data_im_in(978),
            data_im_in(16)=>data_im_in(1042),
            data_im_in(17)=>data_im_in(1106),
            data_im_in(18)=>data_im_in(1170),
            data_im_in(19)=>data_im_in(1234),
            data_im_in(20)=>data_im_in(1298),
            data_im_in(21)=>data_im_in(1362),
            data_im_in(22)=>data_im_in(1426),
            data_im_in(23)=>data_im_in(1490),
            data_im_in(24)=>data_im_in(1554),
            data_im_in(25)=>data_im_in(1618),
            data_im_in(26)=>data_im_in(1682),
            data_im_in(27)=>data_im_in(1746),
            data_im_in(28)=>data_im_in(1810),
            data_im_in(29)=>data_im_in(1874),
            data_im_in(30)=>data_im_in(1938),
            data_im_in(31)=>data_im_in(2002),
            data_re_out=>first_stage_re_out(607 downto 576),
            data_im_out=>first_stage_im_out(607 downto 576)
        );

    ULFFT_PT32_19 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(19),
            data_re_in(1)=>data_re_in(83),
            data_re_in(2)=>data_re_in(147),
            data_re_in(3)=>data_re_in(211),
            data_re_in(4)=>data_re_in(275),
            data_re_in(5)=>data_re_in(339),
            data_re_in(6)=>data_re_in(403),
            data_re_in(7)=>data_re_in(467),
            data_re_in(8)=>data_re_in(531),
            data_re_in(9)=>data_re_in(595),
            data_re_in(10)=>data_re_in(659),
            data_re_in(11)=>data_re_in(723),
            data_re_in(12)=>data_re_in(787),
            data_re_in(13)=>data_re_in(851),
            data_re_in(14)=>data_re_in(915),
            data_re_in(15)=>data_re_in(979),
            data_re_in(16)=>data_re_in(1043),
            data_re_in(17)=>data_re_in(1107),
            data_re_in(18)=>data_re_in(1171),
            data_re_in(19)=>data_re_in(1235),
            data_re_in(20)=>data_re_in(1299),
            data_re_in(21)=>data_re_in(1363),
            data_re_in(22)=>data_re_in(1427),
            data_re_in(23)=>data_re_in(1491),
            data_re_in(24)=>data_re_in(1555),
            data_re_in(25)=>data_re_in(1619),
            data_re_in(26)=>data_re_in(1683),
            data_re_in(27)=>data_re_in(1747),
            data_re_in(28)=>data_re_in(1811),
            data_re_in(29)=>data_re_in(1875),
            data_re_in(30)=>data_re_in(1939),
            data_re_in(31)=>data_re_in(2003),
            data_im_in(0)=>data_im_in(19),
            data_im_in(1)=>data_im_in(83),
            data_im_in(2)=>data_im_in(147),
            data_im_in(3)=>data_im_in(211),
            data_im_in(4)=>data_im_in(275),
            data_im_in(5)=>data_im_in(339),
            data_im_in(6)=>data_im_in(403),
            data_im_in(7)=>data_im_in(467),
            data_im_in(8)=>data_im_in(531),
            data_im_in(9)=>data_im_in(595),
            data_im_in(10)=>data_im_in(659),
            data_im_in(11)=>data_im_in(723),
            data_im_in(12)=>data_im_in(787),
            data_im_in(13)=>data_im_in(851),
            data_im_in(14)=>data_im_in(915),
            data_im_in(15)=>data_im_in(979),
            data_im_in(16)=>data_im_in(1043),
            data_im_in(17)=>data_im_in(1107),
            data_im_in(18)=>data_im_in(1171),
            data_im_in(19)=>data_im_in(1235),
            data_im_in(20)=>data_im_in(1299),
            data_im_in(21)=>data_im_in(1363),
            data_im_in(22)=>data_im_in(1427),
            data_im_in(23)=>data_im_in(1491),
            data_im_in(24)=>data_im_in(1555),
            data_im_in(25)=>data_im_in(1619),
            data_im_in(26)=>data_im_in(1683),
            data_im_in(27)=>data_im_in(1747),
            data_im_in(28)=>data_im_in(1811),
            data_im_in(29)=>data_im_in(1875),
            data_im_in(30)=>data_im_in(1939),
            data_im_in(31)=>data_im_in(2003),
            data_re_out=>first_stage_re_out(639 downto 608),
            data_im_out=>first_stage_im_out(639 downto 608)
        );

    ULFFT_PT32_20 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(20),
            data_re_in(1)=>data_re_in(84),
            data_re_in(2)=>data_re_in(148),
            data_re_in(3)=>data_re_in(212),
            data_re_in(4)=>data_re_in(276),
            data_re_in(5)=>data_re_in(340),
            data_re_in(6)=>data_re_in(404),
            data_re_in(7)=>data_re_in(468),
            data_re_in(8)=>data_re_in(532),
            data_re_in(9)=>data_re_in(596),
            data_re_in(10)=>data_re_in(660),
            data_re_in(11)=>data_re_in(724),
            data_re_in(12)=>data_re_in(788),
            data_re_in(13)=>data_re_in(852),
            data_re_in(14)=>data_re_in(916),
            data_re_in(15)=>data_re_in(980),
            data_re_in(16)=>data_re_in(1044),
            data_re_in(17)=>data_re_in(1108),
            data_re_in(18)=>data_re_in(1172),
            data_re_in(19)=>data_re_in(1236),
            data_re_in(20)=>data_re_in(1300),
            data_re_in(21)=>data_re_in(1364),
            data_re_in(22)=>data_re_in(1428),
            data_re_in(23)=>data_re_in(1492),
            data_re_in(24)=>data_re_in(1556),
            data_re_in(25)=>data_re_in(1620),
            data_re_in(26)=>data_re_in(1684),
            data_re_in(27)=>data_re_in(1748),
            data_re_in(28)=>data_re_in(1812),
            data_re_in(29)=>data_re_in(1876),
            data_re_in(30)=>data_re_in(1940),
            data_re_in(31)=>data_re_in(2004),
            data_im_in(0)=>data_im_in(20),
            data_im_in(1)=>data_im_in(84),
            data_im_in(2)=>data_im_in(148),
            data_im_in(3)=>data_im_in(212),
            data_im_in(4)=>data_im_in(276),
            data_im_in(5)=>data_im_in(340),
            data_im_in(6)=>data_im_in(404),
            data_im_in(7)=>data_im_in(468),
            data_im_in(8)=>data_im_in(532),
            data_im_in(9)=>data_im_in(596),
            data_im_in(10)=>data_im_in(660),
            data_im_in(11)=>data_im_in(724),
            data_im_in(12)=>data_im_in(788),
            data_im_in(13)=>data_im_in(852),
            data_im_in(14)=>data_im_in(916),
            data_im_in(15)=>data_im_in(980),
            data_im_in(16)=>data_im_in(1044),
            data_im_in(17)=>data_im_in(1108),
            data_im_in(18)=>data_im_in(1172),
            data_im_in(19)=>data_im_in(1236),
            data_im_in(20)=>data_im_in(1300),
            data_im_in(21)=>data_im_in(1364),
            data_im_in(22)=>data_im_in(1428),
            data_im_in(23)=>data_im_in(1492),
            data_im_in(24)=>data_im_in(1556),
            data_im_in(25)=>data_im_in(1620),
            data_im_in(26)=>data_im_in(1684),
            data_im_in(27)=>data_im_in(1748),
            data_im_in(28)=>data_im_in(1812),
            data_im_in(29)=>data_im_in(1876),
            data_im_in(30)=>data_im_in(1940),
            data_im_in(31)=>data_im_in(2004),
            data_re_out=>first_stage_re_out(671 downto 640),
            data_im_out=>first_stage_im_out(671 downto 640)
        );

    ULFFT_PT32_21 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(21),
            data_re_in(1)=>data_re_in(85),
            data_re_in(2)=>data_re_in(149),
            data_re_in(3)=>data_re_in(213),
            data_re_in(4)=>data_re_in(277),
            data_re_in(5)=>data_re_in(341),
            data_re_in(6)=>data_re_in(405),
            data_re_in(7)=>data_re_in(469),
            data_re_in(8)=>data_re_in(533),
            data_re_in(9)=>data_re_in(597),
            data_re_in(10)=>data_re_in(661),
            data_re_in(11)=>data_re_in(725),
            data_re_in(12)=>data_re_in(789),
            data_re_in(13)=>data_re_in(853),
            data_re_in(14)=>data_re_in(917),
            data_re_in(15)=>data_re_in(981),
            data_re_in(16)=>data_re_in(1045),
            data_re_in(17)=>data_re_in(1109),
            data_re_in(18)=>data_re_in(1173),
            data_re_in(19)=>data_re_in(1237),
            data_re_in(20)=>data_re_in(1301),
            data_re_in(21)=>data_re_in(1365),
            data_re_in(22)=>data_re_in(1429),
            data_re_in(23)=>data_re_in(1493),
            data_re_in(24)=>data_re_in(1557),
            data_re_in(25)=>data_re_in(1621),
            data_re_in(26)=>data_re_in(1685),
            data_re_in(27)=>data_re_in(1749),
            data_re_in(28)=>data_re_in(1813),
            data_re_in(29)=>data_re_in(1877),
            data_re_in(30)=>data_re_in(1941),
            data_re_in(31)=>data_re_in(2005),
            data_im_in(0)=>data_im_in(21),
            data_im_in(1)=>data_im_in(85),
            data_im_in(2)=>data_im_in(149),
            data_im_in(3)=>data_im_in(213),
            data_im_in(4)=>data_im_in(277),
            data_im_in(5)=>data_im_in(341),
            data_im_in(6)=>data_im_in(405),
            data_im_in(7)=>data_im_in(469),
            data_im_in(8)=>data_im_in(533),
            data_im_in(9)=>data_im_in(597),
            data_im_in(10)=>data_im_in(661),
            data_im_in(11)=>data_im_in(725),
            data_im_in(12)=>data_im_in(789),
            data_im_in(13)=>data_im_in(853),
            data_im_in(14)=>data_im_in(917),
            data_im_in(15)=>data_im_in(981),
            data_im_in(16)=>data_im_in(1045),
            data_im_in(17)=>data_im_in(1109),
            data_im_in(18)=>data_im_in(1173),
            data_im_in(19)=>data_im_in(1237),
            data_im_in(20)=>data_im_in(1301),
            data_im_in(21)=>data_im_in(1365),
            data_im_in(22)=>data_im_in(1429),
            data_im_in(23)=>data_im_in(1493),
            data_im_in(24)=>data_im_in(1557),
            data_im_in(25)=>data_im_in(1621),
            data_im_in(26)=>data_im_in(1685),
            data_im_in(27)=>data_im_in(1749),
            data_im_in(28)=>data_im_in(1813),
            data_im_in(29)=>data_im_in(1877),
            data_im_in(30)=>data_im_in(1941),
            data_im_in(31)=>data_im_in(2005),
            data_re_out=>first_stage_re_out(703 downto 672),
            data_im_out=>first_stage_im_out(703 downto 672)
        );

    ULFFT_PT32_22 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(22),
            data_re_in(1)=>data_re_in(86),
            data_re_in(2)=>data_re_in(150),
            data_re_in(3)=>data_re_in(214),
            data_re_in(4)=>data_re_in(278),
            data_re_in(5)=>data_re_in(342),
            data_re_in(6)=>data_re_in(406),
            data_re_in(7)=>data_re_in(470),
            data_re_in(8)=>data_re_in(534),
            data_re_in(9)=>data_re_in(598),
            data_re_in(10)=>data_re_in(662),
            data_re_in(11)=>data_re_in(726),
            data_re_in(12)=>data_re_in(790),
            data_re_in(13)=>data_re_in(854),
            data_re_in(14)=>data_re_in(918),
            data_re_in(15)=>data_re_in(982),
            data_re_in(16)=>data_re_in(1046),
            data_re_in(17)=>data_re_in(1110),
            data_re_in(18)=>data_re_in(1174),
            data_re_in(19)=>data_re_in(1238),
            data_re_in(20)=>data_re_in(1302),
            data_re_in(21)=>data_re_in(1366),
            data_re_in(22)=>data_re_in(1430),
            data_re_in(23)=>data_re_in(1494),
            data_re_in(24)=>data_re_in(1558),
            data_re_in(25)=>data_re_in(1622),
            data_re_in(26)=>data_re_in(1686),
            data_re_in(27)=>data_re_in(1750),
            data_re_in(28)=>data_re_in(1814),
            data_re_in(29)=>data_re_in(1878),
            data_re_in(30)=>data_re_in(1942),
            data_re_in(31)=>data_re_in(2006),
            data_im_in(0)=>data_im_in(22),
            data_im_in(1)=>data_im_in(86),
            data_im_in(2)=>data_im_in(150),
            data_im_in(3)=>data_im_in(214),
            data_im_in(4)=>data_im_in(278),
            data_im_in(5)=>data_im_in(342),
            data_im_in(6)=>data_im_in(406),
            data_im_in(7)=>data_im_in(470),
            data_im_in(8)=>data_im_in(534),
            data_im_in(9)=>data_im_in(598),
            data_im_in(10)=>data_im_in(662),
            data_im_in(11)=>data_im_in(726),
            data_im_in(12)=>data_im_in(790),
            data_im_in(13)=>data_im_in(854),
            data_im_in(14)=>data_im_in(918),
            data_im_in(15)=>data_im_in(982),
            data_im_in(16)=>data_im_in(1046),
            data_im_in(17)=>data_im_in(1110),
            data_im_in(18)=>data_im_in(1174),
            data_im_in(19)=>data_im_in(1238),
            data_im_in(20)=>data_im_in(1302),
            data_im_in(21)=>data_im_in(1366),
            data_im_in(22)=>data_im_in(1430),
            data_im_in(23)=>data_im_in(1494),
            data_im_in(24)=>data_im_in(1558),
            data_im_in(25)=>data_im_in(1622),
            data_im_in(26)=>data_im_in(1686),
            data_im_in(27)=>data_im_in(1750),
            data_im_in(28)=>data_im_in(1814),
            data_im_in(29)=>data_im_in(1878),
            data_im_in(30)=>data_im_in(1942),
            data_im_in(31)=>data_im_in(2006),
            data_re_out=>first_stage_re_out(735 downto 704),
            data_im_out=>first_stage_im_out(735 downto 704)
        );

    ULFFT_PT32_23 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(23),
            data_re_in(1)=>data_re_in(87),
            data_re_in(2)=>data_re_in(151),
            data_re_in(3)=>data_re_in(215),
            data_re_in(4)=>data_re_in(279),
            data_re_in(5)=>data_re_in(343),
            data_re_in(6)=>data_re_in(407),
            data_re_in(7)=>data_re_in(471),
            data_re_in(8)=>data_re_in(535),
            data_re_in(9)=>data_re_in(599),
            data_re_in(10)=>data_re_in(663),
            data_re_in(11)=>data_re_in(727),
            data_re_in(12)=>data_re_in(791),
            data_re_in(13)=>data_re_in(855),
            data_re_in(14)=>data_re_in(919),
            data_re_in(15)=>data_re_in(983),
            data_re_in(16)=>data_re_in(1047),
            data_re_in(17)=>data_re_in(1111),
            data_re_in(18)=>data_re_in(1175),
            data_re_in(19)=>data_re_in(1239),
            data_re_in(20)=>data_re_in(1303),
            data_re_in(21)=>data_re_in(1367),
            data_re_in(22)=>data_re_in(1431),
            data_re_in(23)=>data_re_in(1495),
            data_re_in(24)=>data_re_in(1559),
            data_re_in(25)=>data_re_in(1623),
            data_re_in(26)=>data_re_in(1687),
            data_re_in(27)=>data_re_in(1751),
            data_re_in(28)=>data_re_in(1815),
            data_re_in(29)=>data_re_in(1879),
            data_re_in(30)=>data_re_in(1943),
            data_re_in(31)=>data_re_in(2007),
            data_im_in(0)=>data_im_in(23),
            data_im_in(1)=>data_im_in(87),
            data_im_in(2)=>data_im_in(151),
            data_im_in(3)=>data_im_in(215),
            data_im_in(4)=>data_im_in(279),
            data_im_in(5)=>data_im_in(343),
            data_im_in(6)=>data_im_in(407),
            data_im_in(7)=>data_im_in(471),
            data_im_in(8)=>data_im_in(535),
            data_im_in(9)=>data_im_in(599),
            data_im_in(10)=>data_im_in(663),
            data_im_in(11)=>data_im_in(727),
            data_im_in(12)=>data_im_in(791),
            data_im_in(13)=>data_im_in(855),
            data_im_in(14)=>data_im_in(919),
            data_im_in(15)=>data_im_in(983),
            data_im_in(16)=>data_im_in(1047),
            data_im_in(17)=>data_im_in(1111),
            data_im_in(18)=>data_im_in(1175),
            data_im_in(19)=>data_im_in(1239),
            data_im_in(20)=>data_im_in(1303),
            data_im_in(21)=>data_im_in(1367),
            data_im_in(22)=>data_im_in(1431),
            data_im_in(23)=>data_im_in(1495),
            data_im_in(24)=>data_im_in(1559),
            data_im_in(25)=>data_im_in(1623),
            data_im_in(26)=>data_im_in(1687),
            data_im_in(27)=>data_im_in(1751),
            data_im_in(28)=>data_im_in(1815),
            data_im_in(29)=>data_im_in(1879),
            data_im_in(30)=>data_im_in(1943),
            data_im_in(31)=>data_im_in(2007),
            data_re_out=>first_stage_re_out(767 downto 736),
            data_im_out=>first_stage_im_out(767 downto 736)
        );

    ULFFT_PT32_24 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(24),
            data_re_in(1)=>data_re_in(88),
            data_re_in(2)=>data_re_in(152),
            data_re_in(3)=>data_re_in(216),
            data_re_in(4)=>data_re_in(280),
            data_re_in(5)=>data_re_in(344),
            data_re_in(6)=>data_re_in(408),
            data_re_in(7)=>data_re_in(472),
            data_re_in(8)=>data_re_in(536),
            data_re_in(9)=>data_re_in(600),
            data_re_in(10)=>data_re_in(664),
            data_re_in(11)=>data_re_in(728),
            data_re_in(12)=>data_re_in(792),
            data_re_in(13)=>data_re_in(856),
            data_re_in(14)=>data_re_in(920),
            data_re_in(15)=>data_re_in(984),
            data_re_in(16)=>data_re_in(1048),
            data_re_in(17)=>data_re_in(1112),
            data_re_in(18)=>data_re_in(1176),
            data_re_in(19)=>data_re_in(1240),
            data_re_in(20)=>data_re_in(1304),
            data_re_in(21)=>data_re_in(1368),
            data_re_in(22)=>data_re_in(1432),
            data_re_in(23)=>data_re_in(1496),
            data_re_in(24)=>data_re_in(1560),
            data_re_in(25)=>data_re_in(1624),
            data_re_in(26)=>data_re_in(1688),
            data_re_in(27)=>data_re_in(1752),
            data_re_in(28)=>data_re_in(1816),
            data_re_in(29)=>data_re_in(1880),
            data_re_in(30)=>data_re_in(1944),
            data_re_in(31)=>data_re_in(2008),
            data_im_in(0)=>data_im_in(24),
            data_im_in(1)=>data_im_in(88),
            data_im_in(2)=>data_im_in(152),
            data_im_in(3)=>data_im_in(216),
            data_im_in(4)=>data_im_in(280),
            data_im_in(5)=>data_im_in(344),
            data_im_in(6)=>data_im_in(408),
            data_im_in(7)=>data_im_in(472),
            data_im_in(8)=>data_im_in(536),
            data_im_in(9)=>data_im_in(600),
            data_im_in(10)=>data_im_in(664),
            data_im_in(11)=>data_im_in(728),
            data_im_in(12)=>data_im_in(792),
            data_im_in(13)=>data_im_in(856),
            data_im_in(14)=>data_im_in(920),
            data_im_in(15)=>data_im_in(984),
            data_im_in(16)=>data_im_in(1048),
            data_im_in(17)=>data_im_in(1112),
            data_im_in(18)=>data_im_in(1176),
            data_im_in(19)=>data_im_in(1240),
            data_im_in(20)=>data_im_in(1304),
            data_im_in(21)=>data_im_in(1368),
            data_im_in(22)=>data_im_in(1432),
            data_im_in(23)=>data_im_in(1496),
            data_im_in(24)=>data_im_in(1560),
            data_im_in(25)=>data_im_in(1624),
            data_im_in(26)=>data_im_in(1688),
            data_im_in(27)=>data_im_in(1752),
            data_im_in(28)=>data_im_in(1816),
            data_im_in(29)=>data_im_in(1880),
            data_im_in(30)=>data_im_in(1944),
            data_im_in(31)=>data_im_in(2008),
            data_re_out=>first_stage_re_out(799 downto 768),
            data_im_out=>first_stage_im_out(799 downto 768)
        );

    ULFFT_PT32_25 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(25),
            data_re_in(1)=>data_re_in(89),
            data_re_in(2)=>data_re_in(153),
            data_re_in(3)=>data_re_in(217),
            data_re_in(4)=>data_re_in(281),
            data_re_in(5)=>data_re_in(345),
            data_re_in(6)=>data_re_in(409),
            data_re_in(7)=>data_re_in(473),
            data_re_in(8)=>data_re_in(537),
            data_re_in(9)=>data_re_in(601),
            data_re_in(10)=>data_re_in(665),
            data_re_in(11)=>data_re_in(729),
            data_re_in(12)=>data_re_in(793),
            data_re_in(13)=>data_re_in(857),
            data_re_in(14)=>data_re_in(921),
            data_re_in(15)=>data_re_in(985),
            data_re_in(16)=>data_re_in(1049),
            data_re_in(17)=>data_re_in(1113),
            data_re_in(18)=>data_re_in(1177),
            data_re_in(19)=>data_re_in(1241),
            data_re_in(20)=>data_re_in(1305),
            data_re_in(21)=>data_re_in(1369),
            data_re_in(22)=>data_re_in(1433),
            data_re_in(23)=>data_re_in(1497),
            data_re_in(24)=>data_re_in(1561),
            data_re_in(25)=>data_re_in(1625),
            data_re_in(26)=>data_re_in(1689),
            data_re_in(27)=>data_re_in(1753),
            data_re_in(28)=>data_re_in(1817),
            data_re_in(29)=>data_re_in(1881),
            data_re_in(30)=>data_re_in(1945),
            data_re_in(31)=>data_re_in(2009),
            data_im_in(0)=>data_im_in(25),
            data_im_in(1)=>data_im_in(89),
            data_im_in(2)=>data_im_in(153),
            data_im_in(3)=>data_im_in(217),
            data_im_in(4)=>data_im_in(281),
            data_im_in(5)=>data_im_in(345),
            data_im_in(6)=>data_im_in(409),
            data_im_in(7)=>data_im_in(473),
            data_im_in(8)=>data_im_in(537),
            data_im_in(9)=>data_im_in(601),
            data_im_in(10)=>data_im_in(665),
            data_im_in(11)=>data_im_in(729),
            data_im_in(12)=>data_im_in(793),
            data_im_in(13)=>data_im_in(857),
            data_im_in(14)=>data_im_in(921),
            data_im_in(15)=>data_im_in(985),
            data_im_in(16)=>data_im_in(1049),
            data_im_in(17)=>data_im_in(1113),
            data_im_in(18)=>data_im_in(1177),
            data_im_in(19)=>data_im_in(1241),
            data_im_in(20)=>data_im_in(1305),
            data_im_in(21)=>data_im_in(1369),
            data_im_in(22)=>data_im_in(1433),
            data_im_in(23)=>data_im_in(1497),
            data_im_in(24)=>data_im_in(1561),
            data_im_in(25)=>data_im_in(1625),
            data_im_in(26)=>data_im_in(1689),
            data_im_in(27)=>data_im_in(1753),
            data_im_in(28)=>data_im_in(1817),
            data_im_in(29)=>data_im_in(1881),
            data_im_in(30)=>data_im_in(1945),
            data_im_in(31)=>data_im_in(2009),
            data_re_out=>first_stage_re_out(831 downto 800),
            data_im_out=>first_stage_im_out(831 downto 800)
        );

    ULFFT_PT32_26 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(26),
            data_re_in(1)=>data_re_in(90),
            data_re_in(2)=>data_re_in(154),
            data_re_in(3)=>data_re_in(218),
            data_re_in(4)=>data_re_in(282),
            data_re_in(5)=>data_re_in(346),
            data_re_in(6)=>data_re_in(410),
            data_re_in(7)=>data_re_in(474),
            data_re_in(8)=>data_re_in(538),
            data_re_in(9)=>data_re_in(602),
            data_re_in(10)=>data_re_in(666),
            data_re_in(11)=>data_re_in(730),
            data_re_in(12)=>data_re_in(794),
            data_re_in(13)=>data_re_in(858),
            data_re_in(14)=>data_re_in(922),
            data_re_in(15)=>data_re_in(986),
            data_re_in(16)=>data_re_in(1050),
            data_re_in(17)=>data_re_in(1114),
            data_re_in(18)=>data_re_in(1178),
            data_re_in(19)=>data_re_in(1242),
            data_re_in(20)=>data_re_in(1306),
            data_re_in(21)=>data_re_in(1370),
            data_re_in(22)=>data_re_in(1434),
            data_re_in(23)=>data_re_in(1498),
            data_re_in(24)=>data_re_in(1562),
            data_re_in(25)=>data_re_in(1626),
            data_re_in(26)=>data_re_in(1690),
            data_re_in(27)=>data_re_in(1754),
            data_re_in(28)=>data_re_in(1818),
            data_re_in(29)=>data_re_in(1882),
            data_re_in(30)=>data_re_in(1946),
            data_re_in(31)=>data_re_in(2010),
            data_im_in(0)=>data_im_in(26),
            data_im_in(1)=>data_im_in(90),
            data_im_in(2)=>data_im_in(154),
            data_im_in(3)=>data_im_in(218),
            data_im_in(4)=>data_im_in(282),
            data_im_in(5)=>data_im_in(346),
            data_im_in(6)=>data_im_in(410),
            data_im_in(7)=>data_im_in(474),
            data_im_in(8)=>data_im_in(538),
            data_im_in(9)=>data_im_in(602),
            data_im_in(10)=>data_im_in(666),
            data_im_in(11)=>data_im_in(730),
            data_im_in(12)=>data_im_in(794),
            data_im_in(13)=>data_im_in(858),
            data_im_in(14)=>data_im_in(922),
            data_im_in(15)=>data_im_in(986),
            data_im_in(16)=>data_im_in(1050),
            data_im_in(17)=>data_im_in(1114),
            data_im_in(18)=>data_im_in(1178),
            data_im_in(19)=>data_im_in(1242),
            data_im_in(20)=>data_im_in(1306),
            data_im_in(21)=>data_im_in(1370),
            data_im_in(22)=>data_im_in(1434),
            data_im_in(23)=>data_im_in(1498),
            data_im_in(24)=>data_im_in(1562),
            data_im_in(25)=>data_im_in(1626),
            data_im_in(26)=>data_im_in(1690),
            data_im_in(27)=>data_im_in(1754),
            data_im_in(28)=>data_im_in(1818),
            data_im_in(29)=>data_im_in(1882),
            data_im_in(30)=>data_im_in(1946),
            data_im_in(31)=>data_im_in(2010),
            data_re_out=>first_stage_re_out(863 downto 832),
            data_im_out=>first_stage_im_out(863 downto 832)
        );

    ULFFT_PT32_27 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(27),
            data_re_in(1)=>data_re_in(91),
            data_re_in(2)=>data_re_in(155),
            data_re_in(3)=>data_re_in(219),
            data_re_in(4)=>data_re_in(283),
            data_re_in(5)=>data_re_in(347),
            data_re_in(6)=>data_re_in(411),
            data_re_in(7)=>data_re_in(475),
            data_re_in(8)=>data_re_in(539),
            data_re_in(9)=>data_re_in(603),
            data_re_in(10)=>data_re_in(667),
            data_re_in(11)=>data_re_in(731),
            data_re_in(12)=>data_re_in(795),
            data_re_in(13)=>data_re_in(859),
            data_re_in(14)=>data_re_in(923),
            data_re_in(15)=>data_re_in(987),
            data_re_in(16)=>data_re_in(1051),
            data_re_in(17)=>data_re_in(1115),
            data_re_in(18)=>data_re_in(1179),
            data_re_in(19)=>data_re_in(1243),
            data_re_in(20)=>data_re_in(1307),
            data_re_in(21)=>data_re_in(1371),
            data_re_in(22)=>data_re_in(1435),
            data_re_in(23)=>data_re_in(1499),
            data_re_in(24)=>data_re_in(1563),
            data_re_in(25)=>data_re_in(1627),
            data_re_in(26)=>data_re_in(1691),
            data_re_in(27)=>data_re_in(1755),
            data_re_in(28)=>data_re_in(1819),
            data_re_in(29)=>data_re_in(1883),
            data_re_in(30)=>data_re_in(1947),
            data_re_in(31)=>data_re_in(2011),
            data_im_in(0)=>data_im_in(27),
            data_im_in(1)=>data_im_in(91),
            data_im_in(2)=>data_im_in(155),
            data_im_in(3)=>data_im_in(219),
            data_im_in(4)=>data_im_in(283),
            data_im_in(5)=>data_im_in(347),
            data_im_in(6)=>data_im_in(411),
            data_im_in(7)=>data_im_in(475),
            data_im_in(8)=>data_im_in(539),
            data_im_in(9)=>data_im_in(603),
            data_im_in(10)=>data_im_in(667),
            data_im_in(11)=>data_im_in(731),
            data_im_in(12)=>data_im_in(795),
            data_im_in(13)=>data_im_in(859),
            data_im_in(14)=>data_im_in(923),
            data_im_in(15)=>data_im_in(987),
            data_im_in(16)=>data_im_in(1051),
            data_im_in(17)=>data_im_in(1115),
            data_im_in(18)=>data_im_in(1179),
            data_im_in(19)=>data_im_in(1243),
            data_im_in(20)=>data_im_in(1307),
            data_im_in(21)=>data_im_in(1371),
            data_im_in(22)=>data_im_in(1435),
            data_im_in(23)=>data_im_in(1499),
            data_im_in(24)=>data_im_in(1563),
            data_im_in(25)=>data_im_in(1627),
            data_im_in(26)=>data_im_in(1691),
            data_im_in(27)=>data_im_in(1755),
            data_im_in(28)=>data_im_in(1819),
            data_im_in(29)=>data_im_in(1883),
            data_im_in(30)=>data_im_in(1947),
            data_im_in(31)=>data_im_in(2011),
            data_re_out=>first_stage_re_out(895 downto 864),
            data_im_out=>first_stage_im_out(895 downto 864)
        );

    ULFFT_PT32_28 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(28),
            data_re_in(1)=>data_re_in(92),
            data_re_in(2)=>data_re_in(156),
            data_re_in(3)=>data_re_in(220),
            data_re_in(4)=>data_re_in(284),
            data_re_in(5)=>data_re_in(348),
            data_re_in(6)=>data_re_in(412),
            data_re_in(7)=>data_re_in(476),
            data_re_in(8)=>data_re_in(540),
            data_re_in(9)=>data_re_in(604),
            data_re_in(10)=>data_re_in(668),
            data_re_in(11)=>data_re_in(732),
            data_re_in(12)=>data_re_in(796),
            data_re_in(13)=>data_re_in(860),
            data_re_in(14)=>data_re_in(924),
            data_re_in(15)=>data_re_in(988),
            data_re_in(16)=>data_re_in(1052),
            data_re_in(17)=>data_re_in(1116),
            data_re_in(18)=>data_re_in(1180),
            data_re_in(19)=>data_re_in(1244),
            data_re_in(20)=>data_re_in(1308),
            data_re_in(21)=>data_re_in(1372),
            data_re_in(22)=>data_re_in(1436),
            data_re_in(23)=>data_re_in(1500),
            data_re_in(24)=>data_re_in(1564),
            data_re_in(25)=>data_re_in(1628),
            data_re_in(26)=>data_re_in(1692),
            data_re_in(27)=>data_re_in(1756),
            data_re_in(28)=>data_re_in(1820),
            data_re_in(29)=>data_re_in(1884),
            data_re_in(30)=>data_re_in(1948),
            data_re_in(31)=>data_re_in(2012),
            data_im_in(0)=>data_im_in(28),
            data_im_in(1)=>data_im_in(92),
            data_im_in(2)=>data_im_in(156),
            data_im_in(3)=>data_im_in(220),
            data_im_in(4)=>data_im_in(284),
            data_im_in(5)=>data_im_in(348),
            data_im_in(6)=>data_im_in(412),
            data_im_in(7)=>data_im_in(476),
            data_im_in(8)=>data_im_in(540),
            data_im_in(9)=>data_im_in(604),
            data_im_in(10)=>data_im_in(668),
            data_im_in(11)=>data_im_in(732),
            data_im_in(12)=>data_im_in(796),
            data_im_in(13)=>data_im_in(860),
            data_im_in(14)=>data_im_in(924),
            data_im_in(15)=>data_im_in(988),
            data_im_in(16)=>data_im_in(1052),
            data_im_in(17)=>data_im_in(1116),
            data_im_in(18)=>data_im_in(1180),
            data_im_in(19)=>data_im_in(1244),
            data_im_in(20)=>data_im_in(1308),
            data_im_in(21)=>data_im_in(1372),
            data_im_in(22)=>data_im_in(1436),
            data_im_in(23)=>data_im_in(1500),
            data_im_in(24)=>data_im_in(1564),
            data_im_in(25)=>data_im_in(1628),
            data_im_in(26)=>data_im_in(1692),
            data_im_in(27)=>data_im_in(1756),
            data_im_in(28)=>data_im_in(1820),
            data_im_in(29)=>data_im_in(1884),
            data_im_in(30)=>data_im_in(1948),
            data_im_in(31)=>data_im_in(2012),
            data_re_out=>first_stage_re_out(927 downto 896),
            data_im_out=>first_stage_im_out(927 downto 896)
        );

    ULFFT_PT32_29 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(29),
            data_re_in(1)=>data_re_in(93),
            data_re_in(2)=>data_re_in(157),
            data_re_in(3)=>data_re_in(221),
            data_re_in(4)=>data_re_in(285),
            data_re_in(5)=>data_re_in(349),
            data_re_in(6)=>data_re_in(413),
            data_re_in(7)=>data_re_in(477),
            data_re_in(8)=>data_re_in(541),
            data_re_in(9)=>data_re_in(605),
            data_re_in(10)=>data_re_in(669),
            data_re_in(11)=>data_re_in(733),
            data_re_in(12)=>data_re_in(797),
            data_re_in(13)=>data_re_in(861),
            data_re_in(14)=>data_re_in(925),
            data_re_in(15)=>data_re_in(989),
            data_re_in(16)=>data_re_in(1053),
            data_re_in(17)=>data_re_in(1117),
            data_re_in(18)=>data_re_in(1181),
            data_re_in(19)=>data_re_in(1245),
            data_re_in(20)=>data_re_in(1309),
            data_re_in(21)=>data_re_in(1373),
            data_re_in(22)=>data_re_in(1437),
            data_re_in(23)=>data_re_in(1501),
            data_re_in(24)=>data_re_in(1565),
            data_re_in(25)=>data_re_in(1629),
            data_re_in(26)=>data_re_in(1693),
            data_re_in(27)=>data_re_in(1757),
            data_re_in(28)=>data_re_in(1821),
            data_re_in(29)=>data_re_in(1885),
            data_re_in(30)=>data_re_in(1949),
            data_re_in(31)=>data_re_in(2013),
            data_im_in(0)=>data_im_in(29),
            data_im_in(1)=>data_im_in(93),
            data_im_in(2)=>data_im_in(157),
            data_im_in(3)=>data_im_in(221),
            data_im_in(4)=>data_im_in(285),
            data_im_in(5)=>data_im_in(349),
            data_im_in(6)=>data_im_in(413),
            data_im_in(7)=>data_im_in(477),
            data_im_in(8)=>data_im_in(541),
            data_im_in(9)=>data_im_in(605),
            data_im_in(10)=>data_im_in(669),
            data_im_in(11)=>data_im_in(733),
            data_im_in(12)=>data_im_in(797),
            data_im_in(13)=>data_im_in(861),
            data_im_in(14)=>data_im_in(925),
            data_im_in(15)=>data_im_in(989),
            data_im_in(16)=>data_im_in(1053),
            data_im_in(17)=>data_im_in(1117),
            data_im_in(18)=>data_im_in(1181),
            data_im_in(19)=>data_im_in(1245),
            data_im_in(20)=>data_im_in(1309),
            data_im_in(21)=>data_im_in(1373),
            data_im_in(22)=>data_im_in(1437),
            data_im_in(23)=>data_im_in(1501),
            data_im_in(24)=>data_im_in(1565),
            data_im_in(25)=>data_im_in(1629),
            data_im_in(26)=>data_im_in(1693),
            data_im_in(27)=>data_im_in(1757),
            data_im_in(28)=>data_im_in(1821),
            data_im_in(29)=>data_im_in(1885),
            data_im_in(30)=>data_im_in(1949),
            data_im_in(31)=>data_im_in(2013),
            data_re_out=>first_stage_re_out(959 downto 928),
            data_im_out=>first_stage_im_out(959 downto 928)
        );

    ULFFT_PT32_30 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(30),
            data_re_in(1)=>data_re_in(94),
            data_re_in(2)=>data_re_in(158),
            data_re_in(3)=>data_re_in(222),
            data_re_in(4)=>data_re_in(286),
            data_re_in(5)=>data_re_in(350),
            data_re_in(6)=>data_re_in(414),
            data_re_in(7)=>data_re_in(478),
            data_re_in(8)=>data_re_in(542),
            data_re_in(9)=>data_re_in(606),
            data_re_in(10)=>data_re_in(670),
            data_re_in(11)=>data_re_in(734),
            data_re_in(12)=>data_re_in(798),
            data_re_in(13)=>data_re_in(862),
            data_re_in(14)=>data_re_in(926),
            data_re_in(15)=>data_re_in(990),
            data_re_in(16)=>data_re_in(1054),
            data_re_in(17)=>data_re_in(1118),
            data_re_in(18)=>data_re_in(1182),
            data_re_in(19)=>data_re_in(1246),
            data_re_in(20)=>data_re_in(1310),
            data_re_in(21)=>data_re_in(1374),
            data_re_in(22)=>data_re_in(1438),
            data_re_in(23)=>data_re_in(1502),
            data_re_in(24)=>data_re_in(1566),
            data_re_in(25)=>data_re_in(1630),
            data_re_in(26)=>data_re_in(1694),
            data_re_in(27)=>data_re_in(1758),
            data_re_in(28)=>data_re_in(1822),
            data_re_in(29)=>data_re_in(1886),
            data_re_in(30)=>data_re_in(1950),
            data_re_in(31)=>data_re_in(2014),
            data_im_in(0)=>data_im_in(30),
            data_im_in(1)=>data_im_in(94),
            data_im_in(2)=>data_im_in(158),
            data_im_in(3)=>data_im_in(222),
            data_im_in(4)=>data_im_in(286),
            data_im_in(5)=>data_im_in(350),
            data_im_in(6)=>data_im_in(414),
            data_im_in(7)=>data_im_in(478),
            data_im_in(8)=>data_im_in(542),
            data_im_in(9)=>data_im_in(606),
            data_im_in(10)=>data_im_in(670),
            data_im_in(11)=>data_im_in(734),
            data_im_in(12)=>data_im_in(798),
            data_im_in(13)=>data_im_in(862),
            data_im_in(14)=>data_im_in(926),
            data_im_in(15)=>data_im_in(990),
            data_im_in(16)=>data_im_in(1054),
            data_im_in(17)=>data_im_in(1118),
            data_im_in(18)=>data_im_in(1182),
            data_im_in(19)=>data_im_in(1246),
            data_im_in(20)=>data_im_in(1310),
            data_im_in(21)=>data_im_in(1374),
            data_im_in(22)=>data_im_in(1438),
            data_im_in(23)=>data_im_in(1502),
            data_im_in(24)=>data_im_in(1566),
            data_im_in(25)=>data_im_in(1630),
            data_im_in(26)=>data_im_in(1694),
            data_im_in(27)=>data_im_in(1758),
            data_im_in(28)=>data_im_in(1822),
            data_im_in(29)=>data_im_in(1886),
            data_im_in(30)=>data_im_in(1950),
            data_im_in(31)=>data_im_in(2014),
            data_re_out=>first_stage_re_out(991 downto 960),
            data_im_out=>first_stage_im_out(991 downto 960)
        );

    ULFFT_PT32_31 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(31),
            data_re_in(1)=>data_re_in(95),
            data_re_in(2)=>data_re_in(159),
            data_re_in(3)=>data_re_in(223),
            data_re_in(4)=>data_re_in(287),
            data_re_in(5)=>data_re_in(351),
            data_re_in(6)=>data_re_in(415),
            data_re_in(7)=>data_re_in(479),
            data_re_in(8)=>data_re_in(543),
            data_re_in(9)=>data_re_in(607),
            data_re_in(10)=>data_re_in(671),
            data_re_in(11)=>data_re_in(735),
            data_re_in(12)=>data_re_in(799),
            data_re_in(13)=>data_re_in(863),
            data_re_in(14)=>data_re_in(927),
            data_re_in(15)=>data_re_in(991),
            data_re_in(16)=>data_re_in(1055),
            data_re_in(17)=>data_re_in(1119),
            data_re_in(18)=>data_re_in(1183),
            data_re_in(19)=>data_re_in(1247),
            data_re_in(20)=>data_re_in(1311),
            data_re_in(21)=>data_re_in(1375),
            data_re_in(22)=>data_re_in(1439),
            data_re_in(23)=>data_re_in(1503),
            data_re_in(24)=>data_re_in(1567),
            data_re_in(25)=>data_re_in(1631),
            data_re_in(26)=>data_re_in(1695),
            data_re_in(27)=>data_re_in(1759),
            data_re_in(28)=>data_re_in(1823),
            data_re_in(29)=>data_re_in(1887),
            data_re_in(30)=>data_re_in(1951),
            data_re_in(31)=>data_re_in(2015),
            data_im_in(0)=>data_im_in(31),
            data_im_in(1)=>data_im_in(95),
            data_im_in(2)=>data_im_in(159),
            data_im_in(3)=>data_im_in(223),
            data_im_in(4)=>data_im_in(287),
            data_im_in(5)=>data_im_in(351),
            data_im_in(6)=>data_im_in(415),
            data_im_in(7)=>data_im_in(479),
            data_im_in(8)=>data_im_in(543),
            data_im_in(9)=>data_im_in(607),
            data_im_in(10)=>data_im_in(671),
            data_im_in(11)=>data_im_in(735),
            data_im_in(12)=>data_im_in(799),
            data_im_in(13)=>data_im_in(863),
            data_im_in(14)=>data_im_in(927),
            data_im_in(15)=>data_im_in(991),
            data_im_in(16)=>data_im_in(1055),
            data_im_in(17)=>data_im_in(1119),
            data_im_in(18)=>data_im_in(1183),
            data_im_in(19)=>data_im_in(1247),
            data_im_in(20)=>data_im_in(1311),
            data_im_in(21)=>data_im_in(1375),
            data_im_in(22)=>data_im_in(1439),
            data_im_in(23)=>data_im_in(1503),
            data_im_in(24)=>data_im_in(1567),
            data_im_in(25)=>data_im_in(1631),
            data_im_in(26)=>data_im_in(1695),
            data_im_in(27)=>data_im_in(1759),
            data_im_in(28)=>data_im_in(1823),
            data_im_in(29)=>data_im_in(1887),
            data_im_in(30)=>data_im_in(1951),
            data_im_in(31)=>data_im_in(2015),
            data_re_out=>first_stage_re_out(1023 downto 992),
            data_im_out=>first_stage_im_out(1023 downto 992)
        );

    ULFFT_PT32_32 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(32),
            data_re_in(1)=>data_re_in(96),
            data_re_in(2)=>data_re_in(160),
            data_re_in(3)=>data_re_in(224),
            data_re_in(4)=>data_re_in(288),
            data_re_in(5)=>data_re_in(352),
            data_re_in(6)=>data_re_in(416),
            data_re_in(7)=>data_re_in(480),
            data_re_in(8)=>data_re_in(544),
            data_re_in(9)=>data_re_in(608),
            data_re_in(10)=>data_re_in(672),
            data_re_in(11)=>data_re_in(736),
            data_re_in(12)=>data_re_in(800),
            data_re_in(13)=>data_re_in(864),
            data_re_in(14)=>data_re_in(928),
            data_re_in(15)=>data_re_in(992),
            data_re_in(16)=>data_re_in(1056),
            data_re_in(17)=>data_re_in(1120),
            data_re_in(18)=>data_re_in(1184),
            data_re_in(19)=>data_re_in(1248),
            data_re_in(20)=>data_re_in(1312),
            data_re_in(21)=>data_re_in(1376),
            data_re_in(22)=>data_re_in(1440),
            data_re_in(23)=>data_re_in(1504),
            data_re_in(24)=>data_re_in(1568),
            data_re_in(25)=>data_re_in(1632),
            data_re_in(26)=>data_re_in(1696),
            data_re_in(27)=>data_re_in(1760),
            data_re_in(28)=>data_re_in(1824),
            data_re_in(29)=>data_re_in(1888),
            data_re_in(30)=>data_re_in(1952),
            data_re_in(31)=>data_re_in(2016),
            data_im_in(0)=>data_im_in(32),
            data_im_in(1)=>data_im_in(96),
            data_im_in(2)=>data_im_in(160),
            data_im_in(3)=>data_im_in(224),
            data_im_in(4)=>data_im_in(288),
            data_im_in(5)=>data_im_in(352),
            data_im_in(6)=>data_im_in(416),
            data_im_in(7)=>data_im_in(480),
            data_im_in(8)=>data_im_in(544),
            data_im_in(9)=>data_im_in(608),
            data_im_in(10)=>data_im_in(672),
            data_im_in(11)=>data_im_in(736),
            data_im_in(12)=>data_im_in(800),
            data_im_in(13)=>data_im_in(864),
            data_im_in(14)=>data_im_in(928),
            data_im_in(15)=>data_im_in(992),
            data_im_in(16)=>data_im_in(1056),
            data_im_in(17)=>data_im_in(1120),
            data_im_in(18)=>data_im_in(1184),
            data_im_in(19)=>data_im_in(1248),
            data_im_in(20)=>data_im_in(1312),
            data_im_in(21)=>data_im_in(1376),
            data_im_in(22)=>data_im_in(1440),
            data_im_in(23)=>data_im_in(1504),
            data_im_in(24)=>data_im_in(1568),
            data_im_in(25)=>data_im_in(1632),
            data_im_in(26)=>data_im_in(1696),
            data_im_in(27)=>data_im_in(1760),
            data_im_in(28)=>data_im_in(1824),
            data_im_in(29)=>data_im_in(1888),
            data_im_in(30)=>data_im_in(1952),
            data_im_in(31)=>data_im_in(2016),
            data_re_out=>first_stage_re_out(1055 downto 1024),
            data_im_out=>first_stage_im_out(1055 downto 1024)
        );

    ULFFT_PT32_33 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(33),
            data_re_in(1)=>data_re_in(97),
            data_re_in(2)=>data_re_in(161),
            data_re_in(3)=>data_re_in(225),
            data_re_in(4)=>data_re_in(289),
            data_re_in(5)=>data_re_in(353),
            data_re_in(6)=>data_re_in(417),
            data_re_in(7)=>data_re_in(481),
            data_re_in(8)=>data_re_in(545),
            data_re_in(9)=>data_re_in(609),
            data_re_in(10)=>data_re_in(673),
            data_re_in(11)=>data_re_in(737),
            data_re_in(12)=>data_re_in(801),
            data_re_in(13)=>data_re_in(865),
            data_re_in(14)=>data_re_in(929),
            data_re_in(15)=>data_re_in(993),
            data_re_in(16)=>data_re_in(1057),
            data_re_in(17)=>data_re_in(1121),
            data_re_in(18)=>data_re_in(1185),
            data_re_in(19)=>data_re_in(1249),
            data_re_in(20)=>data_re_in(1313),
            data_re_in(21)=>data_re_in(1377),
            data_re_in(22)=>data_re_in(1441),
            data_re_in(23)=>data_re_in(1505),
            data_re_in(24)=>data_re_in(1569),
            data_re_in(25)=>data_re_in(1633),
            data_re_in(26)=>data_re_in(1697),
            data_re_in(27)=>data_re_in(1761),
            data_re_in(28)=>data_re_in(1825),
            data_re_in(29)=>data_re_in(1889),
            data_re_in(30)=>data_re_in(1953),
            data_re_in(31)=>data_re_in(2017),
            data_im_in(0)=>data_im_in(33),
            data_im_in(1)=>data_im_in(97),
            data_im_in(2)=>data_im_in(161),
            data_im_in(3)=>data_im_in(225),
            data_im_in(4)=>data_im_in(289),
            data_im_in(5)=>data_im_in(353),
            data_im_in(6)=>data_im_in(417),
            data_im_in(7)=>data_im_in(481),
            data_im_in(8)=>data_im_in(545),
            data_im_in(9)=>data_im_in(609),
            data_im_in(10)=>data_im_in(673),
            data_im_in(11)=>data_im_in(737),
            data_im_in(12)=>data_im_in(801),
            data_im_in(13)=>data_im_in(865),
            data_im_in(14)=>data_im_in(929),
            data_im_in(15)=>data_im_in(993),
            data_im_in(16)=>data_im_in(1057),
            data_im_in(17)=>data_im_in(1121),
            data_im_in(18)=>data_im_in(1185),
            data_im_in(19)=>data_im_in(1249),
            data_im_in(20)=>data_im_in(1313),
            data_im_in(21)=>data_im_in(1377),
            data_im_in(22)=>data_im_in(1441),
            data_im_in(23)=>data_im_in(1505),
            data_im_in(24)=>data_im_in(1569),
            data_im_in(25)=>data_im_in(1633),
            data_im_in(26)=>data_im_in(1697),
            data_im_in(27)=>data_im_in(1761),
            data_im_in(28)=>data_im_in(1825),
            data_im_in(29)=>data_im_in(1889),
            data_im_in(30)=>data_im_in(1953),
            data_im_in(31)=>data_im_in(2017),
            data_re_out=>first_stage_re_out(1087 downto 1056),
            data_im_out=>first_stage_im_out(1087 downto 1056)
        );

    ULFFT_PT32_34 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(34),
            data_re_in(1)=>data_re_in(98),
            data_re_in(2)=>data_re_in(162),
            data_re_in(3)=>data_re_in(226),
            data_re_in(4)=>data_re_in(290),
            data_re_in(5)=>data_re_in(354),
            data_re_in(6)=>data_re_in(418),
            data_re_in(7)=>data_re_in(482),
            data_re_in(8)=>data_re_in(546),
            data_re_in(9)=>data_re_in(610),
            data_re_in(10)=>data_re_in(674),
            data_re_in(11)=>data_re_in(738),
            data_re_in(12)=>data_re_in(802),
            data_re_in(13)=>data_re_in(866),
            data_re_in(14)=>data_re_in(930),
            data_re_in(15)=>data_re_in(994),
            data_re_in(16)=>data_re_in(1058),
            data_re_in(17)=>data_re_in(1122),
            data_re_in(18)=>data_re_in(1186),
            data_re_in(19)=>data_re_in(1250),
            data_re_in(20)=>data_re_in(1314),
            data_re_in(21)=>data_re_in(1378),
            data_re_in(22)=>data_re_in(1442),
            data_re_in(23)=>data_re_in(1506),
            data_re_in(24)=>data_re_in(1570),
            data_re_in(25)=>data_re_in(1634),
            data_re_in(26)=>data_re_in(1698),
            data_re_in(27)=>data_re_in(1762),
            data_re_in(28)=>data_re_in(1826),
            data_re_in(29)=>data_re_in(1890),
            data_re_in(30)=>data_re_in(1954),
            data_re_in(31)=>data_re_in(2018),
            data_im_in(0)=>data_im_in(34),
            data_im_in(1)=>data_im_in(98),
            data_im_in(2)=>data_im_in(162),
            data_im_in(3)=>data_im_in(226),
            data_im_in(4)=>data_im_in(290),
            data_im_in(5)=>data_im_in(354),
            data_im_in(6)=>data_im_in(418),
            data_im_in(7)=>data_im_in(482),
            data_im_in(8)=>data_im_in(546),
            data_im_in(9)=>data_im_in(610),
            data_im_in(10)=>data_im_in(674),
            data_im_in(11)=>data_im_in(738),
            data_im_in(12)=>data_im_in(802),
            data_im_in(13)=>data_im_in(866),
            data_im_in(14)=>data_im_in(930),
            data_im_in(15)=>data_im_in(994),
            data_im_in(16)=>data_im_in(1058),
            data_im_in(17)=>data_im_in(1122),
            data_im_in(18)=>data_im_in(1186),
            data_im_in(19)=>data_im_in(1250),
            data_im_in(20)=>data_im_in(1314),
            data_im_in(21)=>data_im_in(1378),
            data_im_in(22)=>data_im_in(1442),
            data_im_in(23)=>data_im_in(1506),
            data_im_in(24)=>data_im_in(1570),
            data_im_in(25)=>data_im_in(1634),
            data_im_in(26)=>data_im_in(1698),
            data_im_in(27)=>data_im_in(1762),
            data_im_in(28)=>data_im_in(1826),
            data_im_in(29)=>data_im_in(1890),
            data_im_in(30)=>data_im_in(1954),
            data_im_in(31)=>data_im_in(2018),
            data_re_out=>first_stage_re_out(1119 downto 1088),
            data_im_out=>first_stage_im_out(1119 downto 1088)
        );

    ULFFT_PT32_35 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(35),
            data_re_in(1)=>data_re_in(99),
            data_re_in(2)=>data_re_in(163),
            data_re_in(3)=>data_re_in(227),
            data_re_in(4)=>data_re_in(291),
            data_re_in(5)=>data_re_in(355),
            data_re_in(6)=>data_re_in(419),
            data_re_in(7)=>data_re_in(483),
            data_re_in(8)=>data_re_in(547),
            data_re_in(9)=>data_re_in(611),
            data_re_in(10)=>data_re_in(675),
            data_re_in(11)=>data_re_in(739),
            data_re_in(12)=>data_re_in(803),
            data_re_in(13)=>data_re_in(867),
            data_re_in(14)=>data_re_in(931),
            data_re_in(15)=>data_re_in(995),
            data_re_in(16)=>data_re_in(1059),
            data_re_in(17)=>data_re_in(1123),
            data_re_in(18)=>data_re_in(1187),
            data_re_in(19)=>data_re_in(1251),
            data_re_in(20)=>data_re_in(1315),
            data_re_in(21)=>data_re_in(1379),
            data_re_in(22)=>data_re_in(1443),
            data_re_in(23)=>data_re_in(1507),
            data_re_in(24)=>data_re_in(1571),
            data_re_in(25)=>data_re_in(1635),
            data_re_in(26)=>data_re_in(1699),
            data_re_in(27)=>data_re_in(1763),
            data_re_in(28)=>data_re_in(1827),
            data_re_in(29)=>data_re_in(1891),
            data_re_in(30)=>data_re_in(1955),
            data_re_in(31)=>data_re_in(2019),
            data_im_in(0)=>data_im_in(35),
            data_im_in(1)=>data_im_in(99),
            data_im_in(2)=>data_im_in(163),
            data_im_in(3)=>data_im_in(227),
            data_im_in(4)=>data_im_in(291),
            data_im_in(5)=>data_im_in(355),
            data_im_in(6)=>data_im_in(419),
            data_im_in(7)=>data_im_in(483),
            data_im_in(8)=>data_im_in(547),
            data_im_in(9)=>data_im_in(611),
            data_im_in(10)=>data_im_in(675),
            data_im_in(11)=>data_im_in(739),
            data_im_in(12)=>data_im_in(803),
            data_im_in(13)=>data_im_in(867),
            data_im_in(14)=>data_im_in(931),
            data_im_in(15)=>data_im_in(995),
            data_im_in(16)=>data_im_in(1059),
            data_im_in(17)=>data_im_in(1123),
            data_im_in(18)=>data_im_in(1187),
            data_im_in(19)=>data_im_in(1251),
            data_im_in(20)=>data_im_in(1315),
            data_im_in(21)=>data_im_in(1379),
            data_im_in(22)=>data_im_in(1443),
            data_im_in(23)=>data_im_in(1507),
            data_im_in(24)=>data_im_in(1571),
            data_im_in(25)=>data_im_in(1635),
            data_im_in(26)=>data_im_in(1699),
            data_im_in(27)=>data_im_in(1763),
            data_im_in(28)=>data_im_in(1827),
            data_im_in(29)=>data_im_in(1891),
            data_im_in(30)=>data_im_in(1955),
            data_im_in(31)=>data_im_in(2019),
            data_re_out=>first_stage_re_out(1151 downto 1120),
            data_im_out=>first_stage_im_out(1151 downto 1120)
        );

    ULFFT_PT32_36 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(36),
            data_re_in(1)=>data_re_in(100),
            data_re_in(2)=>data_re_in(164),
            data_re_in(3)=>data_re_in(228),
            data_re_in(4)=>data_re_in(292),
            data_re_in(5)=>data_re_in(356),
            data_re_in(6)=>data_re_in(420),
            data_re_in(7)=>data_re_in(484),
            data_re_in(8)=>data_re_in(548),
            data_re_in(9)=>data_re_in(612),
            data_re_in(10)=>data_re_in(676),
            data_re_in(11)=>data_re_in(740),
            data_re_in(12)=>data_re_in(804),
            data_re_in(13)=>data_re_in(868),
            data_re_in(14)=>data_re_in(932),
            data_re_in(15)=>data_re_in(996),
            data_re_in(16)=>data_re_in(1060),
            data_re_in(17)=>data_re_in(1124),
            data_re_in(18)=>data_re_in(1188),
            data_re_in(19)=>data_re_in(1252),
            data_re_in(20)=>data_re_in(1316),
            data_re_in(21)=>data_re_in(1380),
            data_re_in(22)=>data_re_in(1444),
            data_re_in(23)=>data_re_in(1508),
            data_re_in(24)=>data_re_in(1572),
            data_re_in(25)=>data_re_in(1636),
            data_re_in(26)=>data_re_in(1700),
            data_re_in(27)=>data_re_in(1764),
            data_re_in(28)=>data_re_in(1828),
            data_re_in(29)=>data_re_in(1892),
            data_re_in(30)=>data_re_in(1956),
            data_re_in(31)=>data_re_in(2020),
            data_im_in(0)=>data_im_in(36),
            data_im_in(1)=>data_im_in(100),
            data_im_in(2)=>data_im_in(164),
            data_im_in(3)=>data_im_in(228),
            data_im_in(4)=>data_im_in(292),
            data_im_in(5)=>data_im_in(356),
            data_im_in(6)=>data_im_in(420),
            data_im_in(7)=>data_im_in(484),
            data_im_in(8)=>data_im_in(548),
            data_im_in(9)=>data_im_in(612),
            data_im_in(10)=>data_im_in(676),
            data_im_in(11)=>data_im_in(740),
            data_im_in(12)=>data_im_in(804),
            data_im_in(13)=>data_im_in(868),
            data_im_in(14)=>data_im_in(932),
            data_im_in(15)=>data_im_in(996),
            data_im_in(16)=>data_im_in(1060),
            data_im_in(17)=>data_im_in(1124),
            data_im_in(18)=>data_im_in(1188),
            data_im_in(19)=>data_im_in(1252),
            data_im_in(20)=>data_im_in(1316),
            data_im_in(21)=>data_im_in(1380),
            data_im_in(22)=>data_im_in(1444),
            data_im_in(23)=>data_im_in(1508),
            data_im_in(24)=>data_im_in(1572),
            data_im_in(25)=>data_im_in(1636),
            data_im_in(26)=>data_im_in(1700),
            data_im_in(27)=>data_im_in(1764),
            data_im_in(28)=>data_im_in(1828),
            data_im_in(29)=>data_im_in(1892),
            data_im_in(30)=>data_im_in(1956),
            data_im_in(31)=>data_im_in(2020),
            data_re_out=>first_stage_re_out(1183 downto 1152),
            data_im_out=>first_stage_im_out(1183 downto 1152)
        );

    ULFFT_PT32_37 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(37),
            data_re_in(1)=>data_re_in(101),
            data_re_in(2)=>data_re_in(165),
            data_re_in(3)=>data_re_in(229),
            data_re_in(4)=>data_re_in(293),
            data_re_in(5)=>data_re_in(357),
            data_re_in(6)=>data_re_in(421),
            data_re_in(7)=>data_re_in(485),
            data_re_in(8)=>data_re_in(549),
            data_re_in(9)=>data_re_in(613),
            data_re_in(10)=>data_re_in(677),
            data_re_in(11)=>data_re_in(741),
            data_re_in(12)=>data_re_in(805),
            data_re_in(13)=>data_re_in(869),
            data_re_in(14)=>data_re_in(933),
            data_re_in(15)=>data_re_in(997),
            data_re_in(16)=>data_re_in(1061),
            data_re_in(17)=>data_re_in(1125),
            data_re_in(18)=>data_re_in(1189),
            data_re_in(19)=>data_re_in(1253),
            data_re_in(20)=>data_re_in(1317),
            data_re_in(21)=>data_re_in(1381),
            data_re_in(22)=>data_re_in(1445),
            data_re_in(23)=>data_re_in(1509),
            data_re_in(24)=>data_re_in(1573),
            data_re_in(25)=>data_re_in(1637),
            data_re_in(26)=>data_re_in(1701),
            data_re_in(27)=>data_re_in(1765),
            data_re_in(28)=>data_re_in(1829),
            data_re_in(29)=>data_re_in(1893),
            data_re_in(30)=>data_re_in(1957),
            data_re_in(31)=>data_re_in(2021),
            data_im_in(0)=>data_im_in(37),
            data_im_in(1)=>data_im_in(101),
            data_im_in(2)=>data_im_in(165),
            data_im_in(3)=>data_im_in(229),
            data_im_in(4)=>data_im_in(293),
            data_im_in(5)=>data_im_in(357),
            data_im_in(6)=>data_im_in(421),
            data_im_in(7)=>data_im_in(485),
            data_im_in(8)=>data_im_in(549),
            data_im_in(9)=>data_im_in(613),
            data_im_in(10)=>data_im_in(677),
            data_im_in(11)=>data_im_in(741),
            data_im_in(12)=>data_im_in(805),
            data_im_in(13)=>data_im_in(869),
            data_im_in(14)=>data_im_in(933),
            data_im_in(15)=>data_im_in(997),
            data_im_in(16)=>data_im_in(1061),
            data_im_in(17)=>data_im_in(1125),
            data_im_in(18)=>data_im_in(1189),
            data_im_in(19)=>data_im_in(1253),
            data_im_in(20)=>data_im_in(1317),
            data_im_in(21)=>data_im_in(1381),
            data_im_in(22)=>data_im_in(1445),
            data_im_in(23)=>data_im_in(1509),
            data_im_in(24)=>data_im_in(1573),
            data_im_in(25)=>data_im_in(1637),
            data_im_in(26)=>data_im_in(1701),
            data_im_in(27)=>data_im_in(1765),
            data_im_in(28)=>data_im_in(1829),
            data_im_in(29)=>data_im_in(1893),
            data_im_in(30)=>data_im_in(1957),
            data_im_in(31)=>data_im_in(2021),
            data_re_out=>first_stage_re_out(1215 downto 1184),
            data_im_out=>first_stage_im_out(1215 downto 1184)
        );

    ULFFT_PT32_38 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(38),
            data_re_in(1)=>data_re_in(102),
            data_re_in(2)=>data_re_in(166),
            data_re_in(3)=>data_re_in(230),
            data_re_in(4)=>data_re_in(294),
            data_re_in(5)=>data_re_in(358),
            data_re_in(6)=>data_re_in(422),
            data_re_in(7)=>data_re_in(486),
            data_re_in(8)=>data_re_in(550),
            data_re_in(9)=>data_re_in(614),
            data_re_in(10)=>data_re_in(678),
            data_re_in(11)=>data_re_in(742),
            data_re_in(12)=>data_re_in(806),
            data_re_in(13)=>data_re_in(870),
            data_re_in(14)=>data_re_in(934),
            data_re_in(15)=>data_re_in(998),
            data_re_in(16)=>data_re_in(1062),
            data_re_in(17)=>data_re_in(1126),
            data_re_in(18)=>data_re_in(1190),
            data_re_in(19)=>data_re_in(1254),
            data_re_in(20)=>data_re_in(1318),
            data_re_in(21)=>data_re_in(1382),
            data_re_in(22)=>data_re_in(1446),
            data_re_in(23)=>data_re_in(1510),
            data_re_in(24)=>data_re_in(1574),
            data_re_in(25)=>data_re_in(1638),
            data_re_in(26)=>data_re_in(1702),
            data_re_in(27)=>data_re_in(1766),
            data_re_in(28)=>data_re_in(1830),
            data_re_in(29)=>data_re_in(1894),
            data_re_in(30)=>data_re_in(1958),
            data_re_in(31)=>data_re_in(2022),
            data_im_in(0)=>data_im_in(38),
            data_im_in(1)=>data_im_in(102),
            data_im_in(2)=>data_im_in(166),
            data_im_in(3)=>data_im_in(230),
            data_im_in(4)=>data_im_in(294),
            data_im_in(5)=>data_im_in(358),
            data_im_in(6)=>data_im_in(422),
            data_im_in(7)=>data_im_in(486),
            data_im_in(8)=>data_im_in(550),
            data_im_in(9)=>data_im_in(614),
            data_im_in(10)=>data_im_in(678),
            data_im_in(11)=>data_im_in(742),
            data_im_in(12)=>data_im_in(806),
            data_im_in(13)=>data_im_in(870),
            data_im_in(14)=>data_im_in(934),
            data_im_in(15)=>data_im_in(998),
            data_im_in(16)=>data_im_in(1062),
            data_im_in(17)=>data_im_in(1126),
            data_im_in(18)=>data_im_in(1190),
            data_im_in(19)=>data_im_in(1254),
            data_im_in(20)=>data_im_in(1318),
            data_im_in(21)=>data_im_in(1382),
            data_im_in(22)=>data_im_in(1446),
            data_im_in(23)=>data_im_in(1510),
            data_im_in(24)=>data_im_in(1574),
            data_im_in(25)=>data_im_in(1638),
            data_im_in(26)=>data_im_in(1702),
            data_im_in(27)=>data_im_in(1766),
            data_im_in(28)=>data_im_in(1830),
            data_im_in(29)=>data_im_in(1894),
            data_im_in(30)=>data_im_in(1958),
            data_im_in(31)=>data_im_in(2022),
            data_re_out=>first_stage_re_out(1247 downto 1216),
            data_im_out=>first_stage_im_out(1247 downto 1216)
        );

    ULFFT_PT32_39 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(39),
            data_re_in(1)=>data_re_in(103),
            data_re_in(2)=>data_re_in(167),
            data_re_in(3)=>data_re_in(231),
            data_re_in(4)=>data_re_in(295),
            data_re_in(5)=>data_re_in(359),
            data_re_in(6)=>data_re_in(423),
            data_re_in(7)=>data_re_in(487),
            data_re_in(8)=>data_re_in(551),
            data_re_in(9)=>data_re_in(615),
            data_re_in(10)=>data_re_in(679),
            data_re_in(11)=>data_re_in(743),
            data_re_in(12)=>data_re_in(807),
            data_re_in(13)=>data_re_in(871),
            data_re_in(14)=>data_re_in(935),
            data_re_in(15)=>data_re_in(999),
            data_re_in(16)=>data_re_in(1063),
            data_re_in(17)=>data_re_in(1127),
            data_re_in(18)=>data_re_in(1191),
            data_re_in(19)=>data_re_in(1255),
            data_re_in(20)=>data_re_in(1319),
            data_re_in(21)=>data_re_in(1383),
            data_re_in(22)=>data_re_in(1447),
            data_re_in(23)=>data_re_in(1511),
            data_re_in(24)=>data_re_in(1575),
            data_re_in(25)=>data_re_in(1639),
            data_re_in(26)=>data_re_in(1703),
            data_re_in(27)=>data_re_in(1767),
            data_re_in(28)=>data_re_in(1831),
            data_re_in(29)=>data_re_in(1895),
            data_re_in(30)=>data_re_in(1959),
            data_re_in(31)=>data_re_in(2023),
            data_im_in(0)=>data_im_in(39),
            data_im_in(1)=>data_im_in(103),
            data_im_in(2)=>data_im_in(167),
            data_im_in(3)=>data_im_in(231),
            data_im_in(4)=>data_im_in(295),
            data_im_in(5)=>data_im_in(359),
            data_im_in(6)=>data_im_in(423),
            data_im_in(7)=>data_im_in(487),
            data_im_in(8)=>data_im_in(551),
            data_im_in(9)=>data_im_in(615),
            data_im_in(10)=>data_im_in(679),
            data_im_in(11)=>data_im_in(743),
            data_im_in(12)=>data_im_in(807),
            data_im_in(13)=>data_im_in(871),
            data_im_in(14)=>data_im_in(935),
            data_im_in(15)=>data_im_in(999),
            data_im_in(16)=>data_im_in(1063),
            data_im_in(17)=>data_im_in(1127),
            data_im_in(18)=>data_im_in(1191),
            data_im_in(19)=>data_im_in(1255),
            data_im_in(20)=>data_im_in(1319),
            data_im_in(21)=>data_im_in(1383),
            data_im_in(22)=>data_im_in(1447),
            data_im_in(23)=>data_im_in(1511),
            data_im_in(24)=>data_im_in(1575),
            data_im_in(25)=>data_im_in(1639),
            data_im_in(26)=>data_im_in(1703),
            data_im_in(27)=>data_im_in(1767),
            data_im_in(28)=>data_im_in(1831),
            data_im_in(29)=>data_im_in(1895),
            data_im_in(30)=>data_im_in(1959),
            data_im_in(31)=>data_im_in(2023),
            data_re_out=>first_stage_re_out(1279 downto 1248),
            data_im_out=>first_stage_im_out(1279 downto 1248)
        );

    ULFFT_PT32_40 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(40),
            data_re_in(1)=>data_re_in(104),
            data_re_in(2)=>data_re_in(168),
            data_re_in(3)=>data_re_in(232),
            data_re_in(4)=>data_re_in(296),
            data_re_in(5)=>data_re_in(360),
            data_re_in(6)=>data_re_in(424),
            data_re_in(7)=>data_re_in(488),
            data_re_in(8)=>data_re_in(552),
            data_re_in(9)=>data_re_in(616),
            data_re_in(10)=>data_re_in(680),
            data_re_in(11)=>data_re_in(744),
            data_re_in(12)=>data_re_in(808),
            data_re_in(13)=>data_re_in(872),
            data_re_in(14)=>data_re_in(936),
            data_re_in(15)=>data_re_in(1000),
            data_re_in(16)=>data_re_in(1064),
            data_re_in(17)=>data_re_in(1128),
            data_re_in(18)=>data_re_in(1192),
            data_re_in(19)=>data_re_in(1256),
            data_re_in(20)=>data_re_in(1320),
            data_re_in(21)=>data_re_in(1384),
            data_re_in(22)=>data_re_in(1448),
            data_re_in(23)=>data_re_in(1512),
            data_re_in(24)=>data_re_in(1576),
            data_re_in(25)=>data_re_in(1640),
            data_re_in(26)=>data_re_in(1704),
            data_re_in(27)=>data_re_in(1768),
            data_re_in(28)=>data_re_in(1832),
            data_re_in(29)=>data_re_in(1896),
            data_re_in(30)=>data_re_in(1960),
            data_re_in(31)=>data_re_in(2024),
            data_im_in(0)=>data_im_in(40),
            data_im_in(1)=>data_im_in(104),
            data_im_in(2)=>data_im_in(168),
            data_im_in(3)=>data_im_in(232),
            data_im_in(4)=>data_im_in(296),
            data_im_in(5)=>data_im_in(360),
            data_im_in(6)=>data_im_in(424),
            data_im_in(7)=>data_im_in(488),
            data_im_in(8)=>data_im_in(552),
            data_im_in(9)=>data_im_in(616),
            data_im_in(10)=>data_im_in(680),
            data_im_in(11)=>data_im_in(744),
            data_im_in(12)=>data_im_in(808),
            data_im_in(13)=>data_im_in(872),
            data_im_in(14)=>data_im_in(936),
            data_im_in(15)=>data_im_in(1000),
            data_im_in(16)=>data_im_in(1064),
            data_im_in(17)=>data_im_in(1128),
            data_im_in(18)=>data_im_in(1192),
            data_im_in(19)=>data_im_in(1256),
            data_im_in(20)=>data_im_in(1320),
            data_im_in(21)=>data_im_in(1384),
            data_im_in(22)=>data_im_in(1448),
            data_im_in(23)=>data_im_in(1512),
            data_im_in(24)=>data_im_in(1576),
            data_im_in(25)=>data_im_in(1640),
            data_im_in(26)=>data_im_in(1704),
            data_im_in(27)=>data_im_in(1768),
            data_im_in(28)=>data_im_in(1832),
            data_im_in(29)=>data_im_in(1896),
            data_im_in(30)=>data_im_in(1960),
            data_im_in(31)=>data_im_in(2024),
            data_re_out=>first_stage_re_out(1311 downto 1280),
            data_im_out=>first_stage_im_out(1311 downto 1280)
        );

    ULFFT_PT32_41 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(41),
            data_re_in(1)=>data_re_in(105),
            data_re_in(2)=>data_re_in(169),
            data_re_in(3)=>data_re_in(233),
            data_re_in(4)=>data_re_in(297),
            data_re_in(5)=>data_re_in(361),
            data_re_in(6)=>data_re_in(425),
            data_re_in(7)=>data_re_in(489),
            data_re_in(8)=>data_re_in(553),
            data_re_in(9)=>data_re_in(617),
            data_re_in(10)=>data_re_in(681),
            data_re_in(11)=>data_re_in(745),
            data_re_in(12)=>data_re_in(809),
            data_re_in(13)=>data_re_in(873),
            data_re_in(14)=>data_re_in(937),
            data_re_in(15)=>data_re_in(1001),
            data_re_in(16)=>data_re_in(1065),
            data_re_in(17)=>data_re_in(1129),
            data_re_in(18)=>data_re_in(1193),
            data_re_in(19)=>data_re_in(1257),
            data_re_in(20)=>data_re_in(1321),
            data_re_in(21)=>data_re_in(1385),
            data_re_in(22)=>data_re_in(1449),
            data_re_in(23)=>data_re_in(1513),
            data_re_in(24)=>data_re_in(1577),
            data_re_in(25)=>data_re_in(1641),
            data_re_in(26)=>data_re_in(1705),
            data_re_in(27)=>data_re_in(1769),
            data_re_in(28)=>data_re_in(1833),
            data_re_in(29)=>data_re_in(1897),
            data_re_in(30)=>data_re_in(1961),
            data_re_in(31)=>data_re_in(2025),
            data_im_in(0)=>data_im_in(41),
            data_im_in(1)=>data_im_in(105),
            data_im_in(2)=>data_im_in(169),
            data_im_in(3)=>data_im_in(233),
            data_im_in(4)=>data_im_in(297),
            data_im_in(5)=>data_im_in(361),
            data_im_in(6)=>data_im_in(425),
            data_im_in(7)=>data_im_in(489),
            data_im_in(8)=>data_im_in(553),
            data_im_in(9)=>data_im_in(617),
            data_im_in(10)=>data_im_in(681),
            data_im_in(11)=>data_im_in(745),
            data_im_in(12)=>data_im_in(809),
            data_im_in(13)=>data_im_in(873),
            data_im_in(14)=>data_im_in(937),
            data_im_in(15)=>data_im_in(1001),
            data_im_in(16)=>data_im_in(1065),
            data_im_in(17)=>data_im_in(1129),
            data_im_in(18)=>data_im_in(1193),
            data_im_in(19)=>data_im_in(1257),
            data_im_in(20)=>data_im_in(1321),
            data_im_in(21)=>data_im_in(1385),
            data_im_in(22)=>data_im_in(1449),
            data_im_in(23)=>data_im_in(1513),
            data_im_in(24)=>data_im_in(1577),
            data_im_in(25)=>data_im_in(1641),
            data_im_in(26)=>data_im_in(1705),
            data_im_in(27)=>data_im_in(1769),
            data_im_in(28)=>data_im_in(1833),
            data_im_in(29)=>data_im_in(1897),
            data_im_in(30)=>data_im_in(1961),
            data_im_in(31)=>data_im_in(2025),
            data_re_out=>first_stage_re_out(1343 downto 1312),
            data_im_out=>first_stage_im_out(1343 downto 1312)
        );

    ULFFT_PT32_42 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(42),
            data_re_in(1)=>data_re_in(106),
            data_re_in(2)=>data_re_in(170),
            data_re_in(3)=>data_re_in(234),
            data_re_in(4)=>data_re_in(298),
            data_re_in(5)=>data_re_in(362),
            data_re_in(6)=>data_re_in(426),
            data_re_in(7)=>data_re_in(490),
            data_re_in(8)=>data_re_in(554),
            data_re_in(9)=>data_re_in(618),
            data_re_in(10)=>data_re_in(682),
            data_re_in(11)=>data_re_in(746),
            data_re_in(12)=>data_re_in(810),
            data_re_in(13)=>data_re_in(874),
            data_re_in(14)=>data_re_in(938),
            data_re_in(15)=>data_re_in(1002),
            data_re_in(16)=>data_re_in(1066),
            data_re_in(17)=>data_re_in(1130),
            data_re_in(18)=>data_re_in(1194),
            data_re_in(19)=>data_re_in(1258),
            data_re_in(20)=>data_re_in(1322),
            data_re_in(21)=>data_re_in(1386),
            data_re_in(22)=>data_re_in(1450),
            data_re_in(23)=>data_re_in(1514),
            data_re_in(24)=>data_re_in(1578),
            data_re_in(25)=>data_re_in(1642),
            data_re_in(26)=>data_re_in(1706),
            data_re_in(27)=>data_re_in(1770),
            data_re_in(28)=>data_re_in(1834),
            data_re_in(29)=>data_re_in(1898),
            data_re_in(30)=>data_re_in(1962),
            data_re_in(31)=>data_re_in(2026),
            data_im_in(0)=>data_im_in(42),
            data_im_in(1)=>data_im_in(106),
            data_im_in(2)=>data_im_in(170),
            data_im_in(3)=>data_im_in(234),
            data_im_in(4)=>data_im_in(298),
            data_im_in(5)=>data_im_in(362),
            data_im_in(6)=>data_im_in(426),
            data_im_in(7)=>data_im_in(490),
            data_im_in(8)=>data_im_in(554),
            data_im_in(9)=>data_im_in(618),
            data_im_in(10)=>data_im_in(682),
            data_im_in(11)=>data_im_in(746),
            data_im_in(12)=>data_im_in(810),
            data_im_in(13)=>data_im_in(874),
            data_im_in(14)=>data_im_in(938),
            data_im_in(15)=>data_im_in(1002),
            data_im_in(16)=>data_im_in(1066),
            data_im_in(17)=>data_im_in(1130),
            data_im_in(18)=>data_im_in(1194),
            data_im_in(19)=>data_im_in(1258),
            data_im_in(20)=>data_im_in(1322),
            data_im_in(21)=>data_im_in(1386),
            data_im_in(22)=>data_im_in(1450),
            data_im_in(23)=>data_im_in(1514),
            data_im_in(24)=>data_im_in(1578),
            data_im_in(25)=>data_im_in(1642),
            data_im_in(26)=>data_im_in(1706),
            data_im_in(27)=>data_im_in(1770),
            data_im_in(28)=>data_im_in(1834),
            data_im_in(29)=>data_im_in(1898),
            data_im_in(30)=>data_im_in(1962),
            data_im_in(31)=>data_im_in(2026),
            data_re_out=>first_stage_re_out(1375 downto 1344),
            data_im_out=>first_stage_im_out(1375 downto 1344)
        );

    ULFFT_PT32_43 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(43),
            data_re_in(1)=>data_re_in(107),
            data_re_in(2)=>data_re_in(171),
            data_re_in(3)=>data_re_in(235),
            data_re_in(4)=>data_re_in(299),
            data_re_in(5)=>data_re_in(363),
            data_re_in(6)=>data_re_in(427),
            data_re_in(7)=>data_re_in(491),
            data_re_in(8)=>data_re_in(555),
            data_re_in(9)=>data_re_in(619),
            data_re_in(10)=>data_re_in(683),
            data_re_in(11)=>data_re_in(747),
            data_re_in(12)=>data_re_in(811),
            data_re_in(13)=>data_re_in(875),
            data_re_in(14)=>data_re_in(939),
            data_re_in(15)=>data_re_in(1003),
            data_re_in(16)=>data_re_in(1067),
            data_re_in(17)=>data_re_in(1131),
            data_re_in(18)=>data_re_in(1195),
            data_re_in(19)=>data_re_in(1259),
            data_re_in(20)=>data_re_in(1323),
            data_re_in(21)=>data_re_in(1387),
            data_re_in(22)=>data_re_in(1451),
            data_re_in(23)=>data_re_in(1515),
            data_re_in(24)=>data_re_in(1579),
            data_re_in(25)=>data_re_in(1643),
            data_re_in(26)=>data_re_in(1707),
            data_re_in(27)=>data_re_in(1771),
            data_re_in(28)=>data_re_in(1835),
            data_re_in(29)=>data_re_in(1899),
            data_re_in(30)=>data_re_in(1963),
            data_re_in(31)=>data_re_in(2027),
            data_im_in(0)=>data_im_in(43),
            data_im_in(1)=>data_im_in(107),
            data_im_in(2)=>data_im_in(171),
            data_im_in(3)=>data_im_in(235),
            data_im_in(4)=>data_im_in(299),
            data_im_in(5)=>data_im_in(363),
            data_im_in(6)=>data_im_in(427),
            data_im_in(7)=>data_im_in(491),
            data_im_in(8)=>data_im_in(555),
            data_im_in(9)=>data_im_in(619),
            data_im_in(10)=>data_im_in(683),
            data_im_in(11)=>data_im_in(747),
            data_im_in(12)=>data_im_in(811),
            data_im_in(13)=>data_im_in(875),
            data_im_in(14)=>data_im_in(939),
            data_im_in(15)=>data_im_in(1003),
            data_im_in(16)=>data_im_in(1067),
            data_im_in(17)=>data_im_in(1131),
            data_im_in(18)=>data_im_in(1195),
            data_im_in(19)=>data_im_in(1259),
            data_im_in(20)=>data_im_in(1323),
            data_im_in(21)=>data_im_in(1387),
            data_im_in(22)=>data_im_in(1451),
            data_im_in(23)=>data_im_in(1515),
            data_im_in(24)=>data_im_in(1579),
            data_im_in(25)=>data_im_in(1643),
            data_im_in(26)=>data_im_in(1707),
            data_im_in(27)=>data_im_in(1771),
            data_im_in(28)=>data_im_in(1835),
            data_im_in(29)=>data_im_in(1899),
            data_im_in(30)=>data_im_in(1963),
            data_im_in(31)=>data_im_in(2027),
            data_re_out=>first_stage_re_out(1407 downto 1376),
            data_im_out=>first_stage_im_out(1407 downto 1376)
        );

    ULFFT_PT32_44 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(44),
            data_re_in(1)=>data_re_in(108),
            data_re_in(2)=>data_re_in(172),
            data_re_in(3)=>data_re_in(236),
            data_re_in(4)=>data_re_in(300),
            data_re_in(5)=>data_re_in(364),
            data_re_in(6)=>data_re_in(428),
            data_re_in(7)=>data_re_in(492),
            data_re_in(8)=>data_re_in(556),
            data_re_in(9)=>data_re_in(620),
            data_re_in(10)=>data_re_in(684),
            data_re_in(11)=>data_re_in(748),
            data_re_in(12)=>data_re_in(812),
            data_re_in(13)=>data_re_in(876),
            data_re_in(14)=>data_re_in(940),
            data_re_in(15)=>data_re_in(1004),
            data_re_in(16)=>data_re_in(1068),
            data_re_in(17)=>data_re_in(1132),
            data_re_in(18)=>data_re_in(1196),
            data_re_in(19)=>data_re_in(1260),
            data_re_in(20)=>data_re_in(1324),
            data_re_in(21)=>data_re_in(1388),
            data_re_in(22)=>data_re_in(1452),
            data_re_in(23)=>data_re_in(1516),
            data_re_in(24)=>data_re_in(1580),
            data_re_in(25)=>data_re_in(1644),
            data_re_in(26)=>data_re_in(1708),
            data_re_in(27)=>data_re_in(1772),
            data_re_in(28)=>data_re_in(1836),
            data_re_in(29)=>data_re_in(1900),
            data_re_in(30)=>data_re_in(1964),
            data_re_in(31)=>data_re_in(2028),
            data_im_in(0)=>data_im_in(44),
            data_im_in(1)=>data_im_in(108),
            data_im_in(2)=>data_im_in(172),
            data_im_in(3)=>data_im_in(236),
            data_im_in(4)=>data_im_in(300),
            data_im_in(5)=>data_im_in(364),
            data_im_in(6)=>data_im_in(428),
            data_im_in(7)=>data_im_in(492),
            data_im_in(8)=>data_im_in(556),
            data_im_in(9)=>data_im_in(620),
            data_im_in(10)=>data_im_in(684),
            data_im_in(11)=>data_im_in(748),
            data_im_in(12)=>data_im_in(812),
            data_im_in(13)=>data_im_in(876),
            data_im_in(14)=>data_im_in(940),
            data_im_in(15)=>data_im_in(1004),
            data_im_in(16)=>data_im_in(1068),
            data_im_in(17)=>data_im_in(1132),
            data_im_in(18)=>data_im_in(1196),
            data_im_in(19)=>data_im_in(1260),
            data_im_in(20)=>data_im_in(1324),
            data_im_in(21)=>data_im_in(1388),
            data_im_in(22)=>data_im_in(1452),
            data_im_in(23)=>data_im_in(1516),
            data_im_in(24)=>data_im_in(1580),
            data_im_in(25)=>data_im_in(1644),
            data_im_in(26)=>data_im_in(1708),
            data_im_in(27)=>data_im_in(1772),
            data_im_in(28)=>data_im_in(1836),
            data_im_in(29)=>data_im_in(1900),
            data_im_in(30)=>data_im_in(1964),
            data_im_in(31)=>data_im_in(2028),
            data_re_out=>first_stage_re_out(1439 downto 1408),
            data_im_out=>first_stage_im_out(1439 downto 1408)
        );

    ULFFT_PT32_45 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(45),
            data_re_in(1)=>data_re_in(109),
            data_re_in(2)=>data_re_in(173),
            data_re_in(3)=>data_re_in(237),
            data_re_in(4)=>data_re_in(301),
            data_re_in(5)=>data_re_in(365),
            data_re_in(6)=>data_re_in(429),
            data_re_in(7)=>data_re_in(493),
            data_re_in(8)=>data_re_in(557),
            data_re_in(9)=>data_re_in(621),
            data_re_in(10)=>data_re_in(685),
            data_re_in(11)=>data_re_in(749),
            data_re_in(12)=>data_re_in(813),
            data_re_in(13)=>data_re_in(877),
            data_re_in(14)=>data_re_in(941),
            data_re_in(15)=>data_re_in(1005),
            data_re_in(16)=>data_re_in(1069),
            data_re_in(17)=>data_re_in(1133),
            data_re_in(18)=>data_re_in(1197),
            data_re_in(19)=>data_re_in(1261),
            data_re_in(20)=>data_re_in(1325),
            data_re_in(21)=>data_re_in(1389),
            data_re_in(22)=>data_re_in(1453),
            data_re_in(23)=>data_re_in(1517),
            data_re_in(24)=>data_re_in(1581),
            data_re_in(25)=>data_re_in(1645),
            data_re_in(26)=>data_re_in(1709),
            data_re_in(27)=>data_re_in(1773),
            data_re_in(28)=>data_re_in(1837),
            data_re_in(29)=>data_re_in(1901),
            data_re_in(30)=>data_re_in(1965),
            data_re_in(31)=>data_re_in(2029),
            data_im_in(0)=>data_im_in(45),
            data_im_in(1)=>data_im_in(109),
            data_im_in(2)=>data_im_in(173),
            data_im_in(3)=>data_im_in(237),
            data_im_in(4)=>data_im_in(301),
            data_im_in(5)=>data_im_in(365),
            data_im_in(6)=>data_im_in(429),
            data_im_in(7)=>data_im_in(493),
            data_im_in(8)=>data_im_in(557),
            data_im_in(9)=>data_im_in(621),
            data_im_in(10)=>data_im_in(685),
            data_im_in(11)=>data_im_in(749),
            data_im_in(12)=>data_im_in(813),
            data_im_in(13)=>data_im_in(877),
            data_im_in(14)=>data_im_in(941),
            data_im_in(15)=>data_im_in(1005),
            data_im_in(16)=>data_im_in(1069),
            data_im_in(17)=>data_im_in(1133),
            data_im_in(18)=>data_im_in(1197),
            data_im_in(19)=>data_im_in(1261),
            data_im_in(20)=>data_im_in(1325),
            data_im_in(21)=>data_im_in(1389),
            data_im_in(22)=>data_im_in(1453),
            data_im_in(23)=>data_im_in(1517),
            data_im_in(24)=>data_im_in(1581),
            data_im_in(25)=>data_im_in(1645),
            data_im_in(26)=>data_im_in(1709),
            data_im_in(27)=>data_im_in(1773),
            data_im_in(28)=>data_im_in(1837),
            data_im_in(29)=>data_im_in(1901),
            data_im_in(30)=>data_im_in(1965),
            data_im_in(31)=>data_im_in(2029),
            data_re_out=>first_stage_re_out(1471 downto 1440),
            data_im_out=>first_stage_im_out(1471 downto 1440)
        );

    ULFFT_PT32_46 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(46),
            data_re_in(1)=>data_re_in(110),
            data_re_in(2)=>data_re_in(174),
            data_re_in(3)=>data_re_in(238),
            data_re_in(4)=>data_re_in(302),
            data_re_in(5)=>data_re_in(366),
            data_re_in(6)=>data_re_in(430),
            data_re_in(7)=>data_re_in(494),
            data_re_in(8)=>data_re_in(558),
            data_re_in(9)=>data_re_in(622),
            data_re_in(10)=>data_re_in(686),
            data_re_in(11)=>data_re_in(750),
            data_re_in(12)=>data_re_in(814),
            data_re_in(13)=>data_re_in(878),
            data_re_in(14)=>data_re_in(942),
            data_re_in(15)=>data_re_in(1006),
            data_re_in(16)=>data_re_in(1070),
            data_re_in(17)=>data_re_in(1134),
            data_re_in(18)=>data_re_in(1198),
            data_re_in(19)=>data_re_in(1262),
            data_re_in(20)=>data_re_in(1326),
            data_re_in(21)=>data_re_in(1390),
            data_re_in(22)=>data_re_in(1454),
            data_re_in(23)=>data_re_in(1518),
            data_re_in(24)=>data_re_in(1582),
            data_re_in(25)=>data_re_in(1646),
            data_re_in(26)=>data_re_in(1710),
            data_re_in(27)=>data_re_in(1774),
            data_re_in(28)=>data_re_in(1838),
            data_re_in(29)=>data_re_in(1902),
            data_re_in(30)=>data_re_in(1966),
            data_re_in(31)=>data_re_in(2030),
            data_im_in(0)=>data_im_in(46),
            data_im_in(1)=>data_im_in(110),
            data_im_in(2)=>data_im_in(174),
            data_im_in(3)=>data_im_in(238),
            data_im_in(4)=>data_im_in(302),
            data_im_in(5)=>data_im_in(366),
            data_im_in(6)=>data_im_in(430),
            data_im_in(7)=>data_im_in(494),
            data_im_in(8)=>data_im_in(558),
            data_im_in(9)=>data_im_in(622),
            data_im_in(10)=>data_im_in(686),
            data_im_in(11)=>data_im_in(750),
            data_im_in(12)=>data_im_in(814),
            data_im_in(13)=>data_im_in(878),
            data_im_in(14)=>data_im_in(942),
            data_im_in(15)=>data_im_in(1006),
            data_im_in(16)=>data_im_in(1070),
            data_im_in(17)=>data_im_in(1134),
            data_im_in(18)=>data_im_in(1198),
            data_im_in(19)=>data_im_in(1262),
            data_im_in(20)=>data_im_in(1326),
            data_im_in(21)=>data_im_in(1390),
            data_im_in(22)=>data_im_in(1454),
            data_im_in(23)=>data_im_in(1518),
            data_im_in(24)=>data_im_in(1582),
            data_im_in(25)=>data_im_in(1646),
            data_im_in(26)=>data_im_in(1710),
            data_im_in(27)=>data_im_in(1774),
            data_im_in(28)=>data_im_in(1838),
            data_im_in(29)=>data_im_in(1902),
            data_im_in(30)=>data_im_in(1966),
            data_im_in(31)=>data_im_in(2030),
            data_re_out=>first_stage_re_out(1503 downto 1472),
            data_im_out=>first_stage_im_out(1503 downto 1472)
        );

    ULFFT_PT32_47 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(47),
            data_re_in(1)=>data_re_in(111),
            data_re_in(2)=>data_re_in(175),
            data_re_in(3)=>data_re_in(239),
            data_re_in(4)=>data_re_in(303),
            data_re_in(5)=>data_re_in(367),
            data_re_in(6)=>data_re_in(431),
            data_re_in(7)=>data_re_in(495),
            data_re_in(8)=>data_re_in(559),
            data_re_in(9)=>data_re_in(623),
            data_re_in(10)=>data_re_in(687),
            data_re_in(11)=>data_re_in(751),
            data_re_in(12)=>data_re_in(815),
            data_re_in(13)=>data_re_in(879),
            data_re_in(14)=>data_re_in(943),
            data_re_in(15)=>data_re_in(1007),
            data_re_in(16)=>data_re_in(1071),
            data_re_in(17)=>data_re_in(1135),
            data_re_in(18)=>data_re_in(1199),
            data_re_in(19)=>data_re_in(1263),
            data_re_in(20)=>data_re_in(1327),
            data_re_in(21)=>data_re_in(1391),
            data_re_in(22)=>data_re_in(1455),
            data_re_in(23)=>data_re_in(1519),
            data_re_in(24)=>data_re_in(1583),
            data_re_in(25)=>data_re_in(1647),
            data_re_in(26)=>data_re_in(1711),
            data_re_in(27)=>data_re_in(1775),
            data_re_in(28)=>data_re_in(1839),
            data_re_in(29)=>data_re_in(1903),
            data_re_in(30)=>data_re_in(1967),
            data_re_in(31)=>data_re_in(2031),
            data_im_in(0)=>data_im_in(47),
            data_im_in(1)=>data_im_in(111),
            data_im_in(2)=>data_im_in(175),
            data_im_in(3)=>data_im_in(239),
            data_im_in(4)=>data_im_in(303),
            data_im_in(5)=>data_im_in(367),
            data_im_in(6)=>data_im_in(431),
            data_im_in(7)=>data_im_in(495),
            data_im_in(8)=>data_im_in(559),
            data_im_in(9)=>data_im_in(623),
            data_im_in(10)=>data_im_in(687),
            data_im_in(11)=>data_im_in(751),
            data_im_in(12)=>data_im_in(815),
            data_im_in(13)=>data_im_in(879),
            data_im_in(14)=>data_im_in(943),
            data_im_in(15)=>data_im_in(1007),
            data_im_in(16)=>data_im_in(1071),
            data_im_in(17)=>data_im_in(1135),
            data_im_in(18)=>data_im_in(1199),
            data_im_in(19)=>data_im_in(1263),
            data_im_in(20)=>data_im_in(1327),
            data_im_in(21)=>data_im_in(1391),
            data_im_in(22)=>data_im_in(1455),
            data_im_in(23)=>data_im_in(1519),
            data_im_in(24)=>data_im_in(1583),
            data_im_in(25)=>data_im_in(1647),
            data_im_in(26)=>data_im_in(1711),
            data_im_in(27)=>data_im_in(1775),
            data_im_in(28)=>data_im_in(1839),
            data_im_in(29)=>data_im_in(1903),
            data_im_in(30)=>data_im_in(1967),
            data_im_in(31)=>data_im_in(2031),
            data_re_out=>first_stage_re_out(1535 downto 1504),
            data_im_out=>first_stage_im_out(1535 downto 1504)
        );

    ULFFT_PT32_48 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(48),
            data_re_in(1)=>data_re_in(112),
            data_re_in(2)=>data_re_in(176),
            data_re_in(3)=>data_re_in(240),
            data_re_in(4)=>data_re_in(304),
            data_re_in(5)=>data_re_in(368),
            data_re_in(6)=>data_re_in(432),
            data_re_in(7)=>data_re_in(496),
            data_re_in(8)=>data_re_in(560),
            data_re_in(9)=>data_re_in(624),
            data_re_in(10)=>data_re_in(688),
            data_re_in(11)=>data_re_in(752),
            data_re_in(12)=>data_re_in(816),
            data_re_in(13)=>data_re_in(880),
            data_re_in(14)=>data_re_in(944),
            data_re_in(15)=>data_re_in(1008),
            data_re_in(16)=>data_re_in(1072),
            data_re_in(17)=>data_re_in(1136),
            data_re_in(18)=>data_re_in(1200),
            data_re_in(19)=>data_re_in(1264),
            data_re_in(20)=>data_re_in(1328),
            data_re_in(21)=>data_re_in(1392),
            data_re_in(22)=>data_re_in(1456),
            data_re_in(23)=>data_re_in(1520),
            data_re_in(24)=>data_re_in(1584),
            data_re_in(25)=>data_re_in(1648),
            data_re_in(26)=>data_re_in(1712),
            data_re_in(27)=>data_re_in(1776),
            data_re_in(28)=>data_re_in(1840),
            data_re_in(29)=>data_re_in(1904),
            data_re_in(30)=>data_re_in(1968),
            data_re_in(31)=>data_re_in(2032),
            data_im_in(0)=>data_im_in(48),
            data_im_in(1)=>data_im_in(112),
            data_im_in(2)=>data_im_in(176),
            data_im_in(3)=>data_im_in(240),
            data_im_in(4)=>data_im_in(304),
            data_im_in(5)=>data_im_in(368),
            data_im_in(6)=>data_im_in(432),
            data_im_in(7)=>data_im_in(496),
            data_im_in(8)=>data_im_in(560),
            data_im_in(9)=>data_im_in(624),
            data_im_in(10)=>data_im_in(688),
            data_im_in(11)=>data_im_in(752),
            data_im_in(12)=>data_im_in(816),
            data_im_in(13)=>data_im_in(880),
            data_im_in(14)=>data_im_in(944),
            data_im_in(15)=>data_im_in(1008),
            data_im_in(16)=>data_im_in(1072),
            data_im_in(17)=>data_im_in(1136),
            data_im_in(18)=>data_im_in(1200),
            data_im_in(19)=>data_im_in(1264),
            data_im_in(20)=>data_im_in(1328),
            data_im_in(21)=>data_im_in(1392),
            data_im_in(22)=>data_im_in(1456),
            data_im_in(23)=>data_im_in(1520),
            data_im_in(24)=>data_im_in(1584),
            data_im_in(25)=>data_im_in(1648),
            data_im_in(26)=>data_im_in(1712),
            data_im_in(27)=>data_im_in(1776),
            data_im_in(28)=>data_im_in(1840),
            data_im_in(29)=>data_im_in(1904),
            data_im_in(30)=>data_im_in(1968),
            data_im_in(31)=>data_im_in(2032),
            data_re_out=>first_stage_re_out(1567 downto 1536),
            data_im_out=>first_stage_im_out(1567 downto 1536)
        );

    ULFFT_PT32_49 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(49),
            data_re_in(1)=>data_re_in(113),
            data_re_in(2)=>data_re_in(177),
            data_re_in(3)=>data_re_in(241),
            data_re_in(4)=>data_re_in(305),
            data_re_in(5)=>data_re_in(369),
            data_re_in(6)=>data_re_in(433),
            data_re_in(7)=>data_re_in(497),
            data_re_in(8)=>data_re_in(561),
            data_re_in(9)=>data_re_in(625),
            data_re_in(10)=>data_re_in(689),
            data_re_in(11)=>data_re_in(753),
            data_re_in(12)=>data_re_in(817),
            data_re_in(13)=>data_re_in(881),
            data_re_in(14)=>data_re_in(945),
            data_re_in(15)=>data_re_in(1009),
            data_re_in(16)=>data_re_in(1073),
            data_re_in(17)=>data_re_in(1137),
            data_re_in(18)=>data_re_in(1201),
            data_re_in(19)=>data_re_in(1265),
            data_re_in(20)=>data_re_in(1329),
            data_re_in(21)=>data_re_in(1393),
            data_re_in(22)=>data_re_in(1457),
            data_re_in(23)=>data_re_in(1521),
            data_re_in(24)=>data_re_in(1585),
            data_re_in(25)=>data_re_in(1649),
            data_re_in(26)=>data_re_in(1713),
            data_re_in(27)=>data_re_in(1777),
            data_re_in(28)=>data_re_in(1841),
            data_re_in(29)=>data_re_in(1905),
            data_re_in(30)=>data_re_in(1969),
            data_re_in(31)=>data_re_in(2033),
            data_im_in(0)=>data_im_in(49),
            data_im_in(1)=>data_im_in(113),
            data_im_in(2)=>data_im_in(177),
            data_im_in(3)=>data_im_in(241),
            data_im_in(4)=>data_im_in(305),
            data_im_in(5)=>data_im_in(369),
            data_im_in(6)=>data_im_in(433),
            data_im_in(7)=>data_im_in(497),
            data_im_in(8)=>data_im_in(561),
            data_im_in(9)=>data_im_in(625),
            data_im_in(10)=>data_im_in(689),
            data_im_in(11)=>data_im_in(753),
            data_im_in(12)=>data_im_in(817),
            data_im_in(13)=>data_im_in(881),
            data_im_in(14)=>data_im_in(945),
            data_im_in(15)=>data_im_in(1009),
            data_im_in(16)=>data_im_in(1073),
            data_im_in(17)=>data_im_in(1137),
            data_im_in(18)=>data_im_in(1201),
            data_im_in(19)=>data_im_in(1265),
            data_im_in(20)=>data_im_in(1329),
            data_im_in(21)=>data_im_in(1393),
            data_im_in(22)=>data_im_in(1457),
            data_im_in(23)=>data_im_in(1521),
            data_im_in(24)=>data_im_in(1585),
            data_im_in(25)=>data_im_in(1649),
            data_im_in(26)=>data_im_in(1713),
            data_im_in(27)=>data_im_in(1777),
            data_im_in(28)=>data_im_in(1841),
            data_im_in(29)=>data_im_in(1905),
            data_im_in(30)=>data_im_in(1969),
            data_im_in(31)=>data_im_in(2033),
            data_re_out=>first_stage_re_out(1599 downto 1568),
            data_im_out=>first_stage_im_out(1599 downto 1568)
        );

    ULFFT_PT32_50 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(50),
            data_re_in(1)=>data_re_in(114),
            data_re_in(2)=>data_re_in(178),
            data_re_in(3)=>data_re_in(242),
            data_re_in(4)=>data_re_in(306),
            data_re_in(5)=>data_re_in(370),
            data_re_in(6)=>data_re_in(434),
            data_re_in(7)=>data_re_in(498),
            data_re_in(8)=>data_re_in(562),
            data_re_in(9)=>data_re_in(626),
            data_re_in(10)=>data_re_in(690),
            data_re_in(11)=>data_re_in(754),
            data_re_in(12)=>data_re_in(818),
            data_re_in(13)=>data_re_in(882),
            data_re_in(14)=>data_re_in(946),
            data_re_in(15)=>data_re_in(1010),
            data_re_in(16)=>data_re_in(1074),
            data_re_in(17)=>data_re_in(1138),
            data_re_in(18)=>data_re_in(1202),
            data_re_in(19)=>data_re_in(1266),
            data_re_in(20)=>data_re_in(1330),
            data_re_in(21)=>data_re_in(1394),
            data_re_in(22)=>data_re_in(1458),
            data_re_in(23)=>data_re_in(1522),
            data_re_in(24)=>data_re_in(1586),
            data_re_in(25)=>data_re_in(1650),
            data_re_in(26)=>data_re_in(1714),
            data_re_in(27)=>data_re_in(1778),
            data_re_in(28)=>data_re_in(1842),
            data_re_in(29)=>data_re_in(1906),
            data_re_in(30)=>data_re_in(1970),
            data_re_in(31)=>data_re_in(2034),
            data_im_in(0)=>data_im_in(50),
            data_im_in(1)=>data_im_in(114),
            data_im_in(2)=>data_im_in(178),
            data_im_in(3)=>data_im_in(242),
            data_im_in(4)=>data_im_in(306),
            data_im_in(5)=>data_im_in(370),
            data_im_in(6)=>data_im_in(434),
            data_im_in(7)=>data_im_in(498),
            data_im_in(8)=>data_im_in(562),
            data_im_in(9)=>data_im_in(626),
            data_im_in(10)=>data_im_in(690),
            data_im_in(11)=>data_im_in(754),
            data_im_in(12)=>data_im_in(818),
            data_im_in(13)=>data_im_in(882),
            data_im_in(14)=>data_im_in(946),
            data_im_in(15)=>data_im_in(1010),
            data_im_in(16)=>data_im_in(1074),
            data_im_in(17)=>data_im_in(1138),
            data_im_in(18)=>data_im_in(1202),
            data_im_in(19)=>data_im_in(1266),
            data_im_in(20)=>data_im_in(1330),
            data_im_in(21)=>data_im_in(1394),
            data_im_in(22)=>data_im_in(1458),
            data_im_in(23)=>data_im_in(1522),
            data_im_in(24)=>data_im_in(1586),
            data_im_in(25)=>data_im_in(1650),
            data_im_in(26)=>data_im_in(1714),
            data_im_in(27)=>data_im_in(1778),
            data_im_in(28)=>data_im_in(1842),
            data_im_in(29)=>data_im_in(1906),
            data_im_in(30)=>data_im_in(1970),
            data_im_in(31)=>data_im_in(2034),
            data_re_out=>first_stage_re_out(1631 downto 1600),
            data_im_out=>first_stage_im_out(1631 downto 1600)
        );

    ULFFT_PT32_51 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(51),
            data_re_in(1)=>data_re_in(115),
            data_re_in(2)=>data_re_in(179),
            data_re_in(3)=>data_re_in(243),
            data_re_in(4)=>data_re_in(307),
            data_re_in(5)=>data_re_in(371),
            data_re_in(6)=>data_re_in(435),
            data_re_in(7)=>data_re_in(499),
            data_re_in(8)=>data_re_in(563),
            data_re_in(9)=>data_re_in(627),
            data_re_in(10)=>data_re_in(691),
            data_re_in(11)=>data_re_in(755),
            data_re_in(12)=>data_re_in(819),
            data_re_in(13)=>data_re_in(883),
            data_re_in(14)=>data_re_in(947),
            data_re_in(15)=>data_re_in(1011),
            data_re_in(16)=>data_re_in(1075),
            data_re_in(17)=>data_re_in(1139),
            data_re_in(18)=>data_re_in(1203),
            data_re_in(19)=>data_re_in(1267),
            data_re_in(20)=>data_re_in(1331),
            data_re_in(21)=>data_re_in(1395),
            data_re_in(22)=>data_re_in(1459),
            data_re_in(23)=>data_re_in(1523),
            data_re_in(24)=>data_re_in(1587),
            data_re_in(25)=>data_re_in(1651),
            data_re_in(26)=>data_re_in(1715),
            data_re_in(27)=>data_re_in(1779),
            data_re_in(28)=>data_re_in(1843),
            data_re_in(29)=>data_re_in(1907),
            data_re_in(30)=>data_re_in(1971),
            data_re_in(31)=>data_re_in(2035),
            data_im_in(0)=>data_im_in(51),
            data_im_in(1)=>data_im_in(115),
            data_im_in(2)=>data_im_in(179),
            data_im_in(3)=>data_im_in(243),
            data_im_in(4)=>data_im_in(307),
            data_im_in(5)=>data_im_in(371),
            data_im_in(6)=>data_im_in(435),
            data_im_in(7)=>data_im_in(499),
            data_im_in(8)=>data_im_in(563),
            data_im_in(9)=>data_im_in(627),
            data_im_in(10)=>data_im_in(691),
            data_im_in(11)=>data_im_in(755),
            data_im_in(12)=>data_im_in(819),
            data_im_in(13)=>data_im_in(883),
            data_im_in(14)=>data_im_in(947),
            data_im_in(15)=>data_im_in(1011),
            data_im_in(16)=>data_im_in(1075),
            data_im_in(17)=>data_im_in(1139),
            data_im_in(18)=>data_im_in(1203),
            data_im_in(19)=>data_im_in(1267),
            data_im_in(20)=>data_im_in(1331),
            data_im_in(21)=>data_im_in(1395),
            data_im_in(22)=>data_im_in(1459),
            data_im_in(23)=>data_im_in(1523),
            data_im_in(24)=>data_im_in(1587),
            data_im_in(25)=>data_im_in(1651),
            data_im_in(26)=>data_im_in(1715),
            data_im_in(27)=>data_im_in(1779),
            data_im_in(28)=>data_im_in(1843),
            data_im_in(29)=>data_im_in(1907),
            data_im_in(30)=>data_im_in(1971),
            data_im_in(31)=>data_im_in(2035),
            data_re_out=>first_stage_re_out(1663 downto 1632),
            data_im_out=>first_stage_im_out(1663 downto 1632)
        );

    ULFFT_PT32_52 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(52),
            data_re_in(1)=>data_re_in(116),
            data_re_in(2)=>data_re_in(180),
            data_re_in(3)=>data_re_in(244),
            data_re_in(4)=>data_re_in(308),
            data_re_in(5)=>data_re_in(372),
            data_re_in(6)=>data_re_in(436),
            data_re_in(7)=>data_re_in(500),
            data_re_in(8)=>data_re_in(564),
            data_re_in(9)=>data_re_in(628),
            data_re_in(10)=>data_re_in(692),
            data_re_in(11)=>data_re_in(756),
            data_re_in(12)=>data_re_in(820),
            data_re_in(13)=>data_re_in(884),
            data_re_in(14)=>data_re_in(948),
            data_re_in(15)=>data_re_in(1012),
            data_re_in(16)=>data_re_in(1076),
            data_re_in(17)=>data_re_in(1140),
            data_re_in(18)=>data_re_in(1204),
            data_re_in(19)=>data_re_in(1268),
            data_re_in(20)=>data_re_in(1332),
            data_re_in(21)=>data_re_in(1396),
            data_re_in(22)=>data_re_in(1460),
            data_re_in(23)=>data_re_in(1524),
            data_re_in(24)=>data_re_in(1588),
            data_re_in(25)=>data_re_in(1652),
            data_re_in(26)=>data_re_in(1716),
            data_re_in(27)=>data_re_in(1780),
            data_re_in(28)=>data_re_in(1844),
            data_re_in(29)=>data_re_in(1908),
            data_re_in(30)=>data_re_in(1972),
            data_re_in(31)=>data_re_in(2036),
            data_im_in(0)=>data_im_in(52),
            data_im_in(1)=>data_im_in(116),
            data_im_in(2)=>data_im_in(180),
            data_im_in(3)=>data_im_in(244),
            data_im_in(4)=>data_im_in(308),
            data_im_in(5)=>data_im_in(372),
            data_im_in(6)=>data_im_in(436),
            data_im_in(7)=>data_im_in(500),
            data_im_in(8)=>data_im_in(564),
            data_im_in(9)=>data_im_in(628),
            data_im_in(10)=>data_im_in(692),
            data_im_in(11)=>data_im_in(756),
            data_im_in(12)=>data_im_in(820),
            data_im_in(13)=>data_im_in(884),
            data_im_in(14)=>data_im_in(948),
            data_im_in(15)=>data_im_in(1012),
            data_im_in(16)=>data_im_in(1076),
            data_im_in(17)=>data_im_in(1140),
            data_im_in(18)=>data_im_in(1204),
            data_im_in(19)=>data_im_in(1268),
            data_im_in(20)=>data_im_in(1332),
            data_im_in(21)=>data_im_in(1396),
            data_im_in(22)=>data_im_in(1460),
            data_im_in(23)=>data_im_in(1524),
            data_im_in(24)=>data_im_in(1588),
            data_im_in(25)=>data_im_in(1652),
            data_im_in(26)=>data_im_in(1716),
            data_im_in(27)=>data_im_in(1780),
            data_im_in(28)=>data_im_in(1844),
            data_im_in(29)=>data_im_in(1908),
            data_im_in(30)=>data_im_in(1972),
            data_im_in(31)=>data_im_in(2036),
            data_re_out=>first_stage_re_out(1695 downto 1664),
            data_im_out=>first_stage_im_out(1695 downto 1664)
        );

    ULFFT_PT32_53 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(53),
            data_re_in(1)=>data_re_in(117),
            data_re_in(2)=>data_re_in(181),
            data_re_in(3)=>data_re_in(245),
            data_re_in(4)=>data_re_in(309),
            data_re_in(5)=>data_re_in(373),
            data_re_in(6)=>data_re_in(437),
            data_re_in(7)=>data_re_in(501),
            data_re_in(8)=>data_re_in(565),
            data_re_in(9)=>data_re_in(629),
            data_re_in(10)=>data_re_in(693),
            data_re_in(11)=>data_re_in(757),
            data_re_in(12)=>data_re_in(821),
            data_re_in(13)=>data_re_in(885),
            data_re_in(14)=>data_re_in(949),
            data_re_in(15)=>data_re_in(1013),
            data_re_in(16)=>data_re_in(1077),
            data_re_in(17)=>data_re_in(1141),
            data_re_in(18)=>data_re_in(1205),
            data_re_in(19)=>data_re_in(1269),
            data_re_in(20)=>data_re_in(1333),
            data_re_in(21)=>data_re_in(1397),
            data_re_in(22)=>data_re_in(1461),
            data_re_in(23)=>data_re_in(1525),
            data_re_in(24)=>data_re_in(1589),
            data_re_in(25)=>data_re_in(1653),
            data_re_in(26)=>data_re_in(1717),
            data_re_in(27)=>data_re_in(1781),
            data_re_in(28)=>data_re_in(1845),
            data_re_in(29)=>data_re_in(1909),
            data_re_in(30)=>data_re_in(1973),
            data_re_in(31)=>data_re_in(2037),
            data_im_in(0)=>data_im_in(53),
            data_im_in(1)=>data_im_in(117),
            data_im_in(2)=>data_im_in(181),
            data_im_in(3)=>data_im_in(245),
            data_im_in(4)=>data_im_in(309),
            data_im_in(5)=>data_im_in(373),
            data_im_in(6)=>data_im_in(437),
            data_im_in(7)=>data_im_in(501),
            data_im_in(8)=>data_im_in(565),
            data_im_in(9)=>data_im_in(629),
            data_im_in(10)=>data_im_in(693),
            data_im_in(11)=>data_im_in(757),
            data_im_in(12)=>data_im_in(821),
            data_im_in(13)=>data_im_in(885),
            data_im_in(14)=>data_im_in(949),
            data_im_in(15)=>data_im_in(1013),
            data_im_in(16)=>data_im_in(1077),
            data_im_in(17)=>data_im_in(1141),
            data_im_in(18)=>data_im_in(1205),
            data_im_in(19)=>data_im_in(1269),
            data_im_in(20)=>data_im_in(1333),
            data_im_in(21)=>data_im_in(1397),
            data_im_in(22)=>data_im_in(1461),
            data_im_in(23)=>data_im_in(1525),
            data_im_in(24)=>data_im_in(1589),
            data_im_in(25)=>data_im_in(1653),
            data_im_in(26)=>data_im_in(1717),
            data_im_in(27)=>data_im_in(1781),
            data_im_in(28)=>data_im_in(1845),
            data_im_in(29)=>data_im_in(1909),
            data_im_in(30)=>data_im_in(1973),
            data_im_in(31)=>data_im_in(2037),
            data_re_out=>first_stage_re_out(1727 downto 1696),
            data_im_out=>first_stage_im_out(1727 downto 1696)
        );

    ULFFT_PT32_54 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(54),
            data_re_in(1)=>data_re_in(118),
            data_re_in(2)=>data_re_in(182),
            data_re_in(3)=>data_re_in(246),
            data_re_in(4)=>data_re_in(310),
            data_re_in(5)=>data_re_in(374),
            data_re_in(6)=>data_re_in(438),
            data_re_in(7)=>data_re_in(502),
            data_re_in(8)=>data_re_in(566),
            data_re_in(9)=>data_re_in(630),
            data_re_in(10)=>data_re_in(694),
            data_re_in(11)=>data_re_in(758),
            data_re_in(12)=>data_re_in(822),
            data_re_in(13)=>data_re_in(886),
            data_re_in(14)=>data_re_in(950),
            data_re_in(15)=>data_re_in(1014),
            data_re_in(16)=>data_re_in(1078),
            data_re_in(17)=>data_re_in(1142),
            data_re_in(18)=>data_re_in(1206),
            data_re_in(19)=>data_re_in(1270),
            data_re_in(20)=>data_re_in(1334),
            data_re_in(21)=>data_re_in(1398),
            data_re_in(22)=>data_re_in(1462),
            data_re_in(23)=>data_re_in(1526),
            data_re_in(24)=>data_re_in(1590),
            data_re_in(25)=>data_re_in(1654),
            data_re_in(26)=>data_re_in(1718),
            data_re_in(27)=>data_re_in(1782),
            data_re_in(28)=>data_re_in(1846),
            data_re_in(29)=>data_re_in(1910),
            data_re_in(30)=>data_re_in(1974),
            data_re_in(31)=>data_re_in(2038),
            data_im_in(0)=>data_im_in(54),
            data_im_in(1)=>data_im_in(118),
            data_im_in(2)=>data_im_in(182),
            data_im_in(3)=>data_im_in(246),
            data_im_in(4)=>data_im_in(310),
            data_im_in(5)=>data_im_in(374),
            data_im_in(6)=>data_im_in(438),
            data_im_in(7)=>data_im_in(502),
            data_im_in(8)=>data_im_in(566),
            data_im_in(9)=>data_im_in(630),
            data_im_in(10)=>data_im_in(694),
            data_im_in(11)=>data_im_in(758),
            data_im_in(12)=>data_im_in(822),
            data_im_in(13)=>data_im_in(886),
            data_im_in(14)=>data_im_in(950),
            data_im_in(15)=>data_im_in(1014),
            data_im_in(16)=>data_im_in(1078),
            data_im_in(17)=>data_im_in(1142),
            data_im_in(18)=>data_im_in(1206),
            data_im_in(19)=>data_im_in(1270),
            data_im_in(20)=>data_im_in(1334),
            data_im_in(21)=>data_im_in(1398),
            data_im_in(22)=>data_im_in(1462),
            data_im_in(23)=>data_im_in(1526),
            data_im_in(24)=>data_im_in(1590),
            data_im_in(25)=>data_im_in(1654),
            data_im_in(26)=>data_im_in(1718),
            data_im_in(27)=>data_im_in(1782),
            data_im_in(28)=>data_im_in(1846),
            data_im_in(29)=>data_im_in(1910),
            data_im_in(30)=>data_im_in(1974),
            data_im_in(31)=>data_im_in(2038),
            data_re_out=>first_stage_re_out(1759 downto 1728),
            data_im_out=>first_stage_im_out(1759 downto 1728)
        );

    ULFFT_PT32_55 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(55),
            data_re_in(1)=>data_re_in(119),
            data_re_in(2)=>data_re_in(183),
            data_re_in(3)=>data_re_in(247),
            data_re_in(4)=>data_re_in(311),
            data_re_in(5)=>data_re_in(375),
            data_re_in(6)=>data_re_in(439),
            data_re_in(7)=>data_re_in(503),
            data_re_in(8)=>data_re_in(567),
            data_re_in(9)=>data_re_in(631),
            data_re_in(10)=>data_re_in(695),
            data_re_in(11)=>data_re_in(759),
            data_re_in(12)=>data_re_in(823),
            data_re_in(13)=>data_re_in(887),
            data_re_in(14)=>data_re_in(951),
            data_re_in(15)=>data_re_in(1015),
            data_re_in(16)=>data_re_in(1079),
            data_re_in(17)=>data_re_in(1143),
            data_re_in(18)=>data_re_in(1207),
            data_re_in(19)=>data_re_in(1271),
            data_re_in(20)=>data_re_in(1335),
            data_re_in(21)=>data_re_in(1399),
            data_re_in(22)=>data_re_in(1463),
            data_re_in(23)=>data_re_in(1527),
            data_re_in(24)=>data_re_in(1591),
            data_re_in(25)=>data_re_in(1655),
            data_re_in(26)=>data_re_in(1719),
            data_re_in(27)=>data_re_in(1783),
            data_re_in(28)=>data_re_in(1847),
            data_re_in(29)=>data_re_in(1911),
            data_re_in(30)=>data_re_in(1975),
            data_re_in(31)=>data_re_in(2039),
            data_im_in(0)=>data_im_in(55),
            data_im_in(1)=>data_im_in(119),
            data_im_in(2)=>data_im_in(183),
            data_im_in(3)=>data_im_in(247),
            data_im_in(4)=>data_im_in(311),
            data_im_in(5)=>data_im_in(375),
            data_im_in(6)=>data_im_in(439),
            data_im_in(7)=>data_im_in(503),
            data_im_in(8)=>data_im_in(567),
            data_im_in(9)=>data_im_in(631),
            data_im_in(10)=>data_im_in(695),
            data_im_in(11)=>data_im_in(759),
            data_im_in(12)=>data_im_in(823),
            data_im_in(13)=>data_im_in(887),
            data_im_in(14)=>data_im_in(951),
            data_im_in(15)=>data_im_in(1015),
            data_im_in(16)=>data_im_in(1079),
            data_im_in(17)=>data_im_in(1143),
            data_im_in(18)=>data_im_in(1207),
            data_im_in(19)=>data_im_in(1271),
            data_im_in(20)=>data_im_in(1335),
            data_im_in(21)=>data_im_in(1399),
            data_im_in(22)=>data_im_in(1463),
            data_im_in(23)=>data_im_in(1527),
            data_im_in(24)=>data_im_in(1591),
            data_im_in(25)=>data_im_in(1655),
            data_im_in(26)=>data_im_in(1719),
            data_im_in(27)=>data_im_in(1783),
            data_im_in(28)=>data_im_in(1847),
            data_im_in(29)=>data_im_in(1911),
            data_im_in(30)=>data_im_in(1975),
            data_im_in(31)=>data_im_in(2039),
            data_re_out=>first_stage_re_out(1791 downto 1760),
            data_im_out=>first_stage_im_out(1791 downto 1760)
        );

    ULFFT_PT32_56 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(56),
            data_re_in(1)=>data_re_in(120),
            data_re_in(2)=>data_re_in(184),
            data_re_in(3)=>data_re_in(248),
            data_re_in(4)=>data_re_in(312),
            data_re_in(5)=>data_re_in(376),
            data_re_in(6)=>data_re_in(440),
            data_re_in(7)=>data_re_in(504),
            data_re_in(8)=>data_re_in(568),
            data_re_in(9)=>data_re_in(632),
            data_re_in(10)=>data_re_in(696),
            data_re_in(11)=>data_re_in(760),
            data_re_in(12)=>data_re_in(824),
            data_re_in(13)=>data_re_in(888),
            data_re_in(14)=>data_re_in(952),
            data_re_in(15)=>data_re_in(1016),
            data_re_in(16)=>data_re_in(1080),
            data_re_in(17)=>data_re_in(1144),
            data_re_in(18)=>data_re_in(1208),
            data_re_in(19)=>data_re_in(1272),
            data_re_in(20)=>data_re_in(1336),
            data_re_in(21)=>data_re_in(1400),
            data_re_in(22)=>data_re_in(1464),
            data_re_in(23)=>data_re_in(1528),
            data_re_in(24)=>data_re_in(1592),
            data_re_in(25)=>data_re_in(1656),
            data_re_in(26)=>data_re_in(1720),
            data_re_in(27)=>data_re_in(1784),
            data_re_in(28)=>data_re_in(1848),
            data_re_in(29)=>data_re_in(1912),
            data_re_in(30)=>data_re_in(1976),
            data_re_in(31)=>data_re_in(2040),
            data_im_in(0)=>data_im_in(56),
            data_im_in(1)=>data_im_in(120),
            data_im_in(2)=>data_im_in(184),
            data_im_in(3)=>data_im_in(248),
            data_im_in(4)=>data_im_in(312),
            data_im_in(5)=>data_im_in(376),
            data_im_in(6)=>data_im_in(440),
            data_im_in(7)=>data_im_in(504),
            data_im_in(8)=>data_im_in(568),
            data_im_in(9)=>data_im_in(632),
            data_im_in(10)=>data_im_in(696),
            data_im_in(11)=>data_im_in(760),
            data_im_in(12)=>data_im_in(824),
            data_im_in(13)=>data_im_in(888),
            data_im_in(14)=>data_im_in(952),
            data_im_in(15)=>data_im_in(1016),
            data_im_in(16)=>data_im_in(1080),
            data_im_in(17)=>data_im_in(1144),
            data_im_in(18)=>data_im_in(1208),
            data_im_in(19)=>data_im_in(1272),
            data_im_in(20)=>data_im_in(1336),
            data_im_in(21)=>data_im_in(1400),
            data_im_in(22)=>data_im_in(1464),
            data_im_in(23)=>data_im_in(1528),
            data_im_in(24)=>data_im_in(1592),
            data_im_in(25)=>data_im_in(1656),
            data_im_in(26)=>data_im_in(1720),
            data_im_in(27)=>data_im_in(1784),
            data_im_in(28)=>data_im_in(1848),
            data_im_in(29)=>data_im_in(1912),
            data_im_in(30)=>data_im_in(1976),
            data_im_in(31)=>data_im_in(2040),
            data_re_out=>first_stage_re_out(1823 downto 1792),
            data_im_out=>first_stage_im_out(1823 downto 1792)
        );

    ULFFT_PT32_57 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(57),
            data_re_in(1)=>data_re_in(121),
            data_re_in(2)=>data_re_in(185),
            data_re_in(3)=>data_re_in(249),
            data_re_in(4)=>data_re_in(313),
            data_re_in(5)=>data_re_in(377),
            data_re_in(6)=>data_re_in(441),
            data_re_in(7)=>data_re_in(505),
            data_re_in(8)=>data_re_in(569),
            data_re_in(9)=>data_re_in(633),
            data_re_in(10)=>data_re_in(697),
            data_re_in(11)=>data_re_in(761),
            data_re_in(12)=>data_re_in(825),
            data_re_in(13)=>data_re_in(889),
            data_re_in(14)=>data_re_in(953),
            data_re_in(15)=>data_re_in(1017),
            data_re_in(16)=>data_re_in(1081),
            data_re_in(17)=>data_re_in(1145),
            data_re_in(18)=>data_re_in(1209),
            data_re_in(19)=>data_re_in(1273),
            data_re_in(20)=>data_re_in(1337),
            data_re_in(21)=>data_re_in(1401),
            data_re_in(22)=>data_re_in(1465),
            data_re_in(23)=>data_re_in(1529),
            data_re_in(24)=>data_re_in(1593),
            data_re_in(25)=>data_re_in(1657),
            data_re_in(26)=>data_re_in(1721),
            data_re_in(27)=>data_re_in(1785),
            data_re_in(28)=>data_re_in(1849),
            data_re_in(29)=>data_re_in(1913),
            data_re_in(30)=>data_re_in(1977),
            data_re_in(31)=>data_re_in(2041),
            data_im_in(0)=>data_im_in(57),
            data_im_in(1)=>data_im_in(121),
            data_im_in(2)=>data_im_in(185),
            data_im_in(3)=>data_im_in(249),
            data_im_in(4)=>data_im_in(313),
            data_im_in(5)=>data_im_in(377),
            data_im_in(6)=>data_im_in(441),
            data_im_in(7)=>data_im_in(505),
            data_im_in(8)=>data_im_in(569),
            data_im_in(9)=>data_im_in(633),
            data_im_in(10)=>data_im_in(697),
            data_im_in(11)=>data_im_in(761),
            data_im_in(12)=>data_im_in(825),
            data_im_in(13)=>data_im_in(889),
            data_im_in(14)=>data_im_in(953),
            data_im_in(15)=>data_im_in(1017),
            data_im_in(16)=>data_im_in(1081),
            data_im_in(17)=>data_im_in(1145),
            data_im_in(18)=>data_im_in(1209),
            data_im_in(19)=>data_im_in(1273),
            data_im_in(20)=>data_im_in(1337),
            data_im_in(21)=>data_im_in(1401),
            data_im_in(22)=>data_im_in(1465),
            data_im_in(23)=>data_im_in(1529),
            data_im_in(24)=>data_im_in(1593),
            data_im_in(25)=>data_im_in(1657),
            data_im_in(26)=>data_im_in(1721),
            data_im_in(27)=>data_im_in(1785),
            data_im_in(28)=>data_im_in(1849),
            data_im_in(29)=>data_im_in(1913),
            data_im_in(30)=>data_im_in(1977),
            data_im_in(31)=>data_im_in(2041),
            data_re_out=>first_stage_re_out(1855 downto 1824),
            data_im_out=>first_stage_im_out(1855 downto 1824)
        );

    ULFFT_PT32_58 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(58),
            data_re_in(1)=>data_re_in(122),
            data_re_in(2)=>data_re_in(186),
            data_re_in(3)=>data_re_in(250),
            data_re_in(4)=>data_re_in(314),
            data_re_in(5)=>data_re_in(378),
            data_re_in(6)=>data_re_in(442),
            data_re_in(7)=>data_re_in(506),
            data_re_in(8)=>data_re_in(570),
            data_re_in(9)=>data_re_in(634),
            data_re_in(10)=>data_re_in(698),
            data_re_in(11)=>data_re_in(762),
            data_re_in(12)=>data_re_in(826),
            data_re_in(13)=>data_re_in(890),
            data_re_in(14)=>data_re_in(954),
            data_re_in(15)=>data_re_in(1018),
            data_re_in(16)=>data_re_in(1082),
            data_re_in(17)=>data_re_in(1146),
            data_re_in(18)=>data_re_in(1210),
            data_re_in(19)=>data_re_in(1274),
            data_re_in(20)=>data_re_in(1338),
            data_re_in(21)=>data_re_in(1402),
            data_re_in(22)=>data_re_in(1466),
            data_re_in(23)=>data_re_in(1530),
            data_re_in(24)=>data_re_in(1594),
            data_re_in(25)=>data_re_in(1658),
            data_re_in(26)=>data_re_in(1722),
            data_re_in(27)=>data_re_in(1786),
            data_re_in(28)=>data_re_in(1850),
            data_re_in(29)=>data_re_in(1914),
            data_re_in(30)=>data_re_in(1978),
            data_re_in(31)=>data_re_in(2042),
            data_im_in(0)=>data_im_in(58),
            data_im_in(1)=>data_im_in(122),
            data_im_in(2)=>data_im_in(186),
            data_im_in(3)=>data_im_in(250),
            data_im_in(4)=>data_im_in(314),
            data_im_in(5)=>data_im_in(378),
            data_im_in(6)=>data_im_in(442),
            data_im_in(7)=>data_im_in(506),
            data_im_in(8)=>data_im_in(570),
            data_im_in(9)=>data_im_in(634),
            data_im_in(10)=>data_im_in(698),
            data_im_in(11)=>data_im_in(762),
            data_im_in(12)=>data_im_in(826),
            data_im_in(13)=>data_im_in(890),
            data_im_in(14)=>data_im_in(954),
            data_im_in(15)=>data_im_in(1018),
            data_im_in(16)=>data_im_in(1082),
            data_im_in(17)=>data_im_in(1146),
            data_im_in(18)=>data_im_in(1210),
            data_im_in(19)=>data_im_in(1274),
            data_im_in(20)=>data_im_in(1338),
            data_im_in(21)=>data_im_in(1402),
            data_im_in(22)=>data_im_in(1466),
            data_im_in(23)=>data_im_in(1530),
            data_im_in(24)=>data_im_in(1594),
            data_im_in(25)=>data_im_in(1658),
            data_im_in(26)=>data_im_in(1722),
            data_im_in(27)=>data_im_in(1786),
            data_im_in(28)=>data_im_in(1850),
            data_im_in(29)=>data_im_in(1914),
            data_im_in(30)=>data_im_in(1978),
            data_im_in(31)=>data_im_in(2042),
            data_re_out=>first_stage_re_out(1887 downto 1856),
            data_im_out=>first_stage_im_out(1887 downto 1856)
        );

    ULFFT_PT32_59 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(59),
            data_re_in(1)=>data_re_in(123),
            data_re_in(2)=>data_re_in(187),
            data_re_in(3)=>data_re_in(251),
            data_re_in(4)=>data_re_in(315),
            data_re_in(5)=>data_re_in(379),
            data_re_in(6)=>data_re_in(443),
            data_re_in(7)=>data_re_in(507),
            data_re_in(8)=>data_re_in(571),
            data_re_in(9)=>data_re_in(635),
            data_re_in(10)=>data_re_in(699),
            data_re_in(11)=>data_re_in(763),
            data_re_in(12)=>data_re_in(827),
            data_re_in(13)=>data_re_in(891),
            data_re_in(14)=>data_re_in(955),
            data_re_in(15)=>data_re_in(1019),
            data_re_in(16)=>data_re_in(1083),
            data_re_in(17)=>data_re_in(1147),
            data_re_in(18)=>data_re_in(1211),
            data_re_in(19)=>data_re_in(1275),
            data_re_in(20)=>data_re_in(1339),
            data_re_in(21)=>data_re_in(1403),
            data_re_in(22)=>data_re_in(1467),
            data_re_in(23)=>data_re_in(1531),
            data_re_in(24)=>data_re_in(1595),
            data_re_in(25)=>data_re_in(1659),
            data_re_in(26)=>data_re_in(1723),
            data_re_in(27)=>data_re_in(1787),
            data_re_in(28)=>data_re_in(1851),
            data_re_in(29)=>data_re_in(1915),
            data_re_in(30)=>data_re_in(1979),
            data_re_in(31)=>data_re_in(2043),
            data_im_in(0)=>data_im_in(59),
            data_im_in(1)=>data_im_in(123),
            data_im_in(2)=>data_im_in(187),
            data_im_in(3)=>data_im_in(251),
            data_im_in(4)=>data_im_in(315),
            data_im_in(5)=>data_im_in(379),
            data_im_in(6)=>data_im_in(443),
            data_im_in(7)=>data_im_in(507),
            data_im_in(8)=>data_im_in(571),
            data_im_in(9)=>data_im_in(635),
            data_im_in(10)=>data_im_in(699),
            data_im_in(11)=>data_im_in(763),
            data_im_in(12)=>data_im_in(827),
            data_im_in(13)=>data_im_in(891),
            data_im_in(14)=>data_im_in(955),
            data_im_in(15)=>data_im_in(1019),
            data_im_in(16)=>data_im_in(1083),
            data_im_in(17)=>data_im_in(1147),
            data_im_in(18)=>data_im_in(1211),
            data_im_in(19)=>data_im_in(1275),
            data_im_in(20)=>data_im_in(1339),
            data_im_in(21)=>data_im_in(1403),
            data_im_in(22)=>data_im_in(1467),
            data_im_in(23)=>data_im_in(1531),
            data_im_in(24)=>data_im_in(1595),
            data_im_in(25)=>data_im_in(1659),
            data_im_in(26)=>data_im_in(1723),
            data_im_in(27)=>data_im_in(1787),
            data_im_in(28)=>data_im_in(1851),
            data_im_in(29)=>data_im_in(1915),
            data_im_in(30)=>data_im_in(1979),
            data_im_in(31)=>data_im_in(2043),
            data_re_out=>first_stage_re_out(1919 downto 1888),
            data_im_out=>first_stage_im_out(1919 downto 1888)
        );

    ULFFT_PT32_60 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(60),
            data_re_in(1)=>data_re_in(124),
            data_re_in(2)=>data_re_in(188),
            data_re_in(3)=>data_re_in(252),
            data_re_in(4)=>data_re_in(316),
            data_re_in(5)=>data_re_in(380),
            data_re_in(6)=>data_re_in(444),
            data_re_in(7)=>data_re_in(508),
            data_re_in(8)=>data_re_in(572),
            data_re_in(9)=>data_re_in(636),
            data_re_in(10)=>data_re_in(700),
            data_re_in(11)=>data_re_in(764),
            data_re_in(12)=>data_re_in(828),
            data_re_in(13)=>data_re_in(892),
            data_re_in(14)=>data_re_in(956),
            data_re_in(15)=>data_re_in(1020),
            data_re_in(16)=>data_re_in(1084),
            data_re_in(17)=>data_re_in(1148),
            data_re_in(18)=>data_re_in(1212),
            data_re_in(19)=>data_re_in(1276),
            data_re_in(20)=>data_re_in(1340),
            data_re_in(21)=>data_re_in(1404),
            data_re_in(22)=>data_re_in(1468),
            data_re_in(23)=>data_re_in(1532),
            data_re_in(24)=>data_re_in(1596),
            data_re_in(25)=>data_re_in(1660),
            data_re_in(26)=>data_re_in(1724),
            data_re_in(27)=>data_re_in(1788),
            data_re_in(28)=>data_re_in(1852),
            data_re_in(29)=>data_re_in(1916),
            data_re_in(30)=>data_re_in(1980),
            data_re_in(31)=>data_re_in(2044),
            data_im_in(0)=>data_im_in(60),
            data_im_in(1)=>data_im_in(124),
            data_im_in(2)=>data_im_in(188),
            data_im_in(3)=>data_im_in(252),
            data_im_in(4)=>data_im_in(316),
            data_im_in(5)=>data_im_in(380),
            data_im_in(6)=>data_im_in(444),
            data_im_in(7)=>data_im_in(508),
            data_im_in(8)=>data_im_in(572),
            data_im_in(9)=>data_im_in(636),
            data_im_in(10)=>data_im_in(700),
            data_im_in(11)=>data_im_in(764),
            data_im_in(12)=>data_im_in(828),
            data_im_in(13)=>data_im_in(892),
            data_im_in(14)=>data_im_in(956),
            data_im_in(15)=>data_im_in(1020),
            data_im_in(16)=>data_im_in(1084),
            data_im_in(17)=>data_im_in(1148),
            data_im_in(18)=>data_im_in(1212),
            data_im_in(19)=>data_im_in(1276),
            data_im_in(20)=>data_im_in(1340),
            data_im_in(21)=>data_im_in(1404),
            data_im_in(22)=>data_im_in(1468),
            data_im_in(23)=>data_im_in(1532),
            data_im_in(24)=>data_im_in(1596),
            data_im_in(25)=>data_im_in(1660),
            data_im_in(26)=>data_im_in(1724),
            data_im_in(27)=>data_im_in(1788),
            data_im_in(28)=>data_im_in(1852),
            data_im_in(29)=>data_im_in(1916),
            data_im_in(30)=>data_im_in(1980),
            data_im_in(31)=>data_im_in(2044),
            data_re_out=>first_stage_re_out(1951 downto 1920),
            data_im_out=>first_stage_im_out(1951 downto 1920)
        );

    ULFFT_PT32_61 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(61),
            data_re_in(1)=>data_re_in(125),
            data_re_in(2)=>data_re_in(189),
            data_re_in(3)=>data_re_in(253),
            data_re_in(4)=>data_re_in(317),
            data_re_in(5)=>data_re_in(381),
            data_re_in(6)=>data_re_in(445),
            data_re_in(7)=>data_re_in(509),
            data_re_in(8)=>data_re_in(573),
            data_re_in(9)=>data_re_in(637),
            data_re_in(10)=>data_re_in(701),
            data_re_in(11)=>data_re_in(765),
            data_re_in(12)=>data_re_in(829),
            data_re_in(13)=>data_re_in(893),
            data_re_in(14)=>data_re_in(957),
            data_re_in(15)=>data_re_in(1021),
            data_re_in(16)=>data_re_in(1085),
            data_re_in(17)=>data_re_in(1149),
            data_re_in(18)=>data_re_in(1213),
            data_re_in(19)=>data_re_in(1277),
            data_re_in(20)=>data_re_in(1341),
            data_re_in(21)=>data_re_in(1405),
            data_re_in(22)=>data_re_in(1469),
            data_re_in(23)=>data_re_in(1533),
            data_re_in(24)=>data_re_in(1597),
            data_re_in(25)=>data_re_in(1661),
            data_re_in(26)=>data_re_in(1725),
            data_re_in(27)=>data_re_in(1789),
            data_re_in(28)=>data_re_in(1853),
            data_re_in(29)=>data_re_in(1917),
            data_re_in(30)=>data_re_in(1981),
            data_re_in(31)=>data_re_in(2045),
            data_im_in(0)=>data_im_in(61),
            data_im_in(1)=>data_im_in(125),
            data_im_in(2)=>data_im_in(189),
            data_im_in(3)=>data_im_in(253),
            data_im_in(4)=>data_im_in(317),
            data_im_in(5)=>data_im_in(381),
            data_im_in(6)=>data_im_in(445),
            data_im_in(7)=>data_im_in(509),
            data_im_in(8)=>data_im_in(573),
            data_im_in(9)=>data_im_in(637),
            data_im_in(10)=>data_im_in(701),
            data_im_in(11)=>data_im_in(765),
            data_im_in(12)=>data_im_in(829),
            data_im_in(13)=>data_im_in(893),
            data_im_in(14)=>data_im_in(957),
            data_im_in(15)=>data_im_in(1021),
            data_im_in(16)=>data_im_in(1085),
            data_im_in(17)=>data_im_in(1149),
            data_im_in(18)=>data_im_in(1213),
            data_im_in(19)=>data_im_in(1277),
            data_im_in(20)=>data_im_in(1341),
            data_im_in(21)=>data_im_in(1405),
            data_im_in(22)=>data_im_in(1469),
            data_im_in(23)=>data_im_in(1533),
            data_im_in(24)=>data_im_in(1597),
            data_im_in(25)=>data_im_in(1661),
            data_im_in(26)=>data_im_in(1725),
            data_im_in(27)=>data_im_in(1789),
            data_im_in(28)=>data_im_in(1853),
            data_im_in(29)=>data_im_in(1917),
            data_im_in(30)=>data_im_in(1981),
            data_im_in(31)=>data_im_in(2045),
            data_re_out=>first_stage_re_out(1983 downto 1952),
            data_im_out=>first_stage_im_out(1983 downto 1952)
        );

    ULFFT_PT32_62 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(62),
            data_re_in(1)=>data_re_in(126),
            data_re_in(2)=>data_re_in(190),
            data_re_in(3)=>data_re_in(254),
            data_re_in(4)=>data_re_in(318),
            data_re_in(5)=>data_re_in(382),
            data_re_in(6)=>data_re_in(446),
            data_re_in(7)=>data_re_in(510),
            data_re_in(8)=>data_re_in(574),
            data_re_in(9)=>data_re_in(638),
            data_re_in(10)=>data_re_in(702),
            data_re_in(11)=>data_re_in(766),
            data_re_in(12)=>data_re_in(830),
            data_re_in(13)=>data_re_in(894),
            data_re_in(14)=>data_re_in(958),
            data_re_in(15)=>data_re_in(1022),
            data_re_in(16)=>data_re_in(1086),
            data_re_in(17)=>data_re_in(1150),
            data_re_in(18)=>data_re_in(1214),
            data_re_in(19)=>data_re_in(1278),
            data_re_in(20)=>data_re_in(1342),
            data_re_in(21)=>data_re_in(1406),
            data_re_in(22)=>data_re_in(1470),
            data_re_in(23)=>data_re_in(1534),
            data_re_in(24)=>data_re_in(1598),
            data_re_in(25)=>data_re_in(1662),
            data_re_in(26)=>data_re_in(1726),
            data_re_in(27)=>data_re_in(1790),
            data_re_in(28)=>data_re_in(1854),
            data_re_in(29)=>data_re_in(1918),
            data_re_in(30)=>data_re_in(1982),
            data_re_in(31)=>data_re_in(2046),
            data_im_in(0)=>data_im_in(62),
            data_im_in(1)=>data_im_in(126),
            data_im_in(2)=>data_im_in(190),
            data_im_in(3)=>data_im_in(254),
            data_im_in(4)=>data_im_in(318),
            data_im_in(5)=>data_im_in(382),
            data_im_in(6)=>data_im_in(446),
            data_im_in(7)=>data_im_in(510),
            data_im_in(8)=>data_im_in(574),
            data_im_in(9)=>data_im_in(638),
            data_im_in(10)=>data_im_in(702),
            data_im_in(11)=>data_im_in(766),
            data_im_in(12)=>data_im_in(830),
            data_im_in(13)=>data_im_in(894),
            data_im_in(14)=>data_im_in(958),
            data_im_in(15)=>data_im_in(1022),
            data_im_in(16)=>data_im_in(1086),
            data_im_in(17)=>data_im_in(1150),
            data_im_in(18)=>data_im_in(1214),
            data_im_in(19)=>data_im_in(1278),
            data_im_in(20)=>data_im_in(1342),
            data_im_in(21)=>data_im_in(1406),
            data_im_in(22)=>data_im_in(1470),
            data_im_in(23)=>data_im_in(1534),
            data_im_in(24)=>data_im_in(1598),
            data_im_in(25)=>data_im_in(1662),
            data_im_in(26)=>data_im_in(1726),
            data_im_in(27)=>data_im_in(1790),
            data_im_in(28)=>data_im_in(1854),
            data_im_in(29)=>data_im_in(1918),
            data_im_in(30)=>data_im_in(1982),
            data_im_in(31)=>data_im_in(2046),
            data_re_out=>first_stage_re_out(2015 downto 1984),
            data_im_out=>first_stage_im_out(2015 downto 1984)
        );

    ULFFT_PT32_63 : fft_pt32
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl,
            data_re_in(0)=>data_re_in(63),
            data_re_in(1)=>data_re_in(127),
            data_re_in(2)=>data_re_in(191),
            data_re_in(3)=>data_re_in(255),
            data_re_in(4)=>data_re_in(319),
            data_re_in(5)=>data_re_in(383),
            data_re_in(6)=>data_re_in(447),
            data_re_in(7)=>data_re_in(511),
            data_re_in(8)=>data_re_in(575),
            data_re_in(9)=>data_re_in(639),
            data_re_in(10)=>data_re_in(703),
            data_re_in(11)=>data_re_in(767),
            data_re_in(12)=>data_re_in(831),
            data_re_in(13)=>data_re_in(895),
            data_re_in(14)=>data_re_in(959),
            data_re_in(15)=>data_re_in(1023),
            data_re_in(16)=>data_re_in(1087),
            data_re_in(17)=>data_re_in(1151),
            data_re_in(18)=>data_re_in(1215),
            data_re_in(19)=>data_re_in(1279),
            data_re_in(20)=>data_re_in(1343),
            data_re_in(21)=>data_re_in(1407),
            data_re_in(22)=>data_re_in(1471),
            data_re_in(23)=>data_re_in(1535),
            data_re_in(24)=>data_re_in(1599),
            data_re_in(25)=>data_re_in(1663),
            data_re_in(26)=>data_re_in(1727),
            data_re_in(27)=>data_re_in(1791),
            data_re_in(28)=>data_re_in(1855),
            data_re_in(29)=>data_re_in(1919),
            data_re_in(30)=>data_re_in(1983),
            data_re_in(31)=>data_re_in(2047),
            data_im_in(0)=>data_im_in(63),
            data_im_in(1)=>data_im_in(127),
            data_im_in(2)=>data_im_in(191),
            data_im_in(3)=>data_im_in(255),
            data_im_in(4)=>data_im_in(319),
            data_im_in(5)=>data_im_in(383),
            data_im_in(6)=>data_im_in(447),
            data_im_in(7)=>data_im_in(511),
            data_im_in(8)=>data_im_in(575),
            data_im_in(9)=>data_im_in(639),
            data_im_in(10)=>data_im_in(703),
            data_im_in(11)=>data_im_in(767),
            data_im_in(12)=>data_im_in(831),
            data_im_in(13)=>data_im_in(895),
            data_im_in(14)=>data_im_in(959),
            data_im_in(15)=>data_im_in(1023),
            data_im_in(16)=>data_im_in(1087),
            data_im_in(17)=>data_im_in(1151),
            data_im_in(18)=>data_im_in(1215),
            data_im_in(19)=>data_im_in(1279),
            data_im_in(20)=>data_im_in(1343),
            data_im_in(21)=>data_im_in(1407),
            data_im_in(22)=>data_im_in(1471),
            data_im_in(23)=>data_im_in(1535),
            data_im_in(24)=>data_im_in(1599),
            data_im_in(25)=>data_im_in(1663),
            data_im_in(26)=>data_im_in(1727),
            data_im_in(27)=>data_im_in(1791),
            data_im_in(28)=>data_im_in(1855),
            data_im_in(29)=>data_im_in(1919),
            data_im_in(30)=>data_im_in(1983),
            data_im_in(31)=>data_im_in(2047),
            data_re_out=>first_stage_re_out(2047 downto 2016),
            data_im_out=>first_stage_im_out(2047 downto 2016)
        );


    --- right-hand-side processors
    URFFT_PT64_0 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(0),
            data_re_in(1)=>mul_re_out(32),
            data_re_in(2)=>mul_re_out(64),
            data_re_in(3)=>mul_re_out(96),
            data_re_in(4)=>mul_re_out(128),
            data_re_in(5)=>mul_re_out(160),
            data_re_in(6)=>mul_re_out(192),
            data_re_in(7)=>mul_re_out(224),
            data_re_in(8)=>mul_re_out(256),
            data_re_in(9)=>mul_re_out(288),
            data_re_in(10)=>mul_re_out(320),
            data_re_in(11)=>mul_re_out(352),
            data_re_in(12)=>mul_re_out(384),
            data_re_in(13)=>mul_re_out(416),
            data_re_in(14)=>mul_re_out(448),
            data_re_in(15)=>mul_re_out(480),
            data_re_in(16)=>mul_re_out(512),
            data_re_in(17)=>mul_re_out(544),
            data_re_in(18)=>mul_re_out(576),
            data_re_in(19)=>mul_re_out(608),
            data_re_in(20)=>mul_re_out(640),
            data_re_in(21)=>mul_re_out(672),
            data_re_in(22)=>mul_re_out(704),
            data_re_in(23)=>mul_re_out(736),
            data_re_in(24)=>mul_re_out(768),
            data_re_in(25)=>mul_re_out(800),
            data_re_in(26)=>mul_re_out(832),
            data_re_in(27)=>mul_re_out(864),
            data_re_in(28)=>mul_re_out(896),
            data_re_in(29)=>mul_re_out(928),
            data_re_in(30)=>mul_re_out(960),
            data_re_in(31)=>mul_re_out(992),
            data_re_in(32)=>mul_re_out(1024),
            data_re_in(33)=>mul_re_out(1056),
            data_re_in(34)=>mul_re_out(1088),
            data_re_in(35)=>mul_re_out(1120),
            data_re_in(36)=>mul_re_out(1152),
            data_re_in(37)=>mul_re_out(1184),
            data_re_in(38)=>mul_re_out(1216),
            data_re_in(39)=>mul_re_out(1248),
            data_re_in(40)=>mul_re_out(1280),
            data_re_in(41)=>mul_re_out(1312),
            data_re_in(42)=>mul_re_out(1344),
            data_re_in(43)=>mul_re_out(1376),
            data_re_in(44)=>mul_re_out(1408),
            data_re_in(45)=>mul_re_out(1440),
            data_re_in(46)=>mul_re_out(1472),
            data_re_in(47)=>mul_re_out(1504),
            data_re_in(48)=>mul_re_out(1536),
            data_re_in(49)=>mul_re_out(1568),
            data_re_in(50)=>mul_re_out(1600),
            data_re_in(51)=>mul_re_out(1632),
            data_re_in(52)=>mul_re_out(1664),
            data_re_in(53)=>mul_re_out(1696),
            data_re_in(54)=>mul_re_out(1728),
            data_re_in(55)=>mul_re_out(1760),
            data_re_in(56)=>mul_re_out(1792),
            data_re_in(57)=>mul_re_out(1824),
            data_re_in(58)=>mul_re_out(1856),
            data_re_in(59)=>mul_re_out(1888),
            data_re_in(60)=>mul_re_out(1920),
            data_re_in(61)=>mul_re_out(1952),
            data_re_in(62)=>mul_re_out(1984),
            data_re_in(63)=>mul_re_out(2016),
            data_im_in(0)=>mul_im_out(0),
            data_im_in(1)=>mul_im_out(32),
            data_im_in(2)=>mul_im_out(64),
            data_im_in(3)=>mul_im_out(96),
            data_im_in(4)=>mul_im_out(128),
            data_im_in(5)=>mul_im_out(160),
            data_im_in(6)=>mul_im_out(192),
            data_im_in(7)=>mul_im_out(224),
            data_im_in(8)=>mul_im_out(256),
            data_im_in(9)=>mul_im_out(288),
            data_im_in(10)=>mul_im_out(320),
            data_im_in(11)=>mul_im_out(352),
            data_im_in(12)=>mul_im_out(384),
            data_im_in(13)=>mul_im_out(416),
            data_im_in(14)=>mul_im_out(448),
            data_im_in(15)=>mul_im_out(480),
            data_im_in(16)=>mul_im_out(512),
            data_im_in(17)=>mul_im_out(544),
            data_im_in(18)=>mul_im_out(576),
            data_im_in(19)=>mul_im_out(608),
            data_im_in(20)=>mul_im_out(640),
            data_im_in(21)=>mul_im_out(672),
            data_im_in(22)=>mul_im_out(704),
            data_im_in(23)=>mul_im_out(736),
            data_im_in(24)=>mul_im_out(768),
            data_im_in(25)=>mul_im_out(800),
            data_im_in(26)=>mul_im_out(832),
            data_im_in(27)=>mul_im_out(864),
            data_im_in(28)=>mul_im_out(896),
            data_im_in(29)=>mul_im_out(928),
            data_im_in(30)=>mul_im_out(960),
            data_im_in(31)=>mul_im_out(992),
            data_im_in(32)=>mul_im_out(1024),
            data_im_in(33)=>mul_im_out(1056),
            data_im_in(34)=>mul_im_out(1088),
            data_im_in(35)=>mul_im_out(1120),
            data_im_in(36)=>mul_im_out(1152),
            data_im_in(37)=>mul_im_out(1184),
            data_im_in(38)=>mul_im_out(1216),
            data_im_in(39)=>mul_im_out(1248),
            data_im_in(40)=>mul_im_out(1280),
            data_im_in(41)=>mul_im_out(1312),
            data_im_in(42)=>mul_im_out(1344),
            data_im_in(43)=>mul_im_out(1376),
            data_im_in(44)=>mul_im_out(1408),
            data_im_in(45)=>mul_im_out(1440),
            data_im_in(46)=>mul_im_out(1472),
            data_im_in(47)=>mul_im_out(1504),
            data_im_in(48)=>mul_im_out(1536),
            data_im_in(49)=>mul_im_out(1568),
            data_im_in(50)=>mul_im_out(1600),
            data_im_in(51)=>mul_im_out(1632),
            data_im_in(52)=>mul_im_out(1664),
            data_im_in(53)=>mul_im_out(1696),
            data_im_in(54)=>mul_im_out(1728),
            data_im_in(55)=>mul_im_out(1760),
            data_im_in(56)=>mul_im_out(1792),
            data_im_in(57)=>mul_im_out(1824),
            data_im_in(58)=>mul_im_out(1856),
            data_im_in(59)=>mul_im_out(1888),
            data_im_in(60)=>mul_im_out(1920),
            data_im_in(61)=>mul_im_out(1952),
            data_im_in(62)=>mul_im_out(1984),
            data_im_in(63)=>mul_im_out(2016),
            data_re_out(0)=>data_re_out(0),
            data_re_out(1)=>data_re_out(32),
            data_re_out(2)=>data_re_out(64),
            data_re_out(3)=>data_re_out(96),
            data_re_out(4)=>data_re_out(128),
            data_re_out(5)=>data_re_out(160),
            data_re_out(6)=>data_re_out(192),
            data_re_out(7)=>data_re_out(224),
            data_re_out(8)=>data_re_out(256),
            data_re_out(9)=>data_re_out(288),
            data_re_out(10)=>data_re_out(320),
            data_re_out(11)=>data_re_out(352),
            data_re_out(12)=>data_re_out(384),
            data_re_out(13)=>data_re_out(416),
            data_re_out(14)=>data_re_out(448),
            data_re_out(15)=>data_re_out(480),
            data_re_out(16)=>data_re_out(512),
            data_re_out(17)=>data_re_out(544),
            data_re_out(18)=>data_re_out(576),
            data_re_out(19)=>data_re_out(608),
            data_re_out(20)=>data_re_out(640),
            data_re_out(21)=>data_re_out(672),
            data_re_out(22)=>data_re_out(704),
            data_re_out(23)=>data_re_out(736),
            data_re_out(24)=>data_re_out(768),
            data_re_out(25)=>data_re_out(800),
            data_re_out(26)=>data_re_out(832),
            data_re_out(27)=>data_re_out(864),
            data_re_out(28)=>data_re_out(896),
            data_re_out(29)=>data_re_out(928),
            data_re_out(30)=>data_re_out(960),
            data_re_out(31)=>data_re_out(992),
            data_re_out(32)=>data_re_out(1024),
            data_re_out(33)=>data_re_out(1056),
            data_re_out(34)=>data_re_out(1088),
            data_re_out(35)=>data_re_out(1120),
            data_re_out(36)=>data_re_out(1152),
            data_re_out(37)=>data_re_out(1184),
            data_re_out(38)=>data_re_out(1216),
            data_re_out(39)=>data_re_out(1248),
            data_re_out(40)=>data_re_out(1280),
            data_re_out(41)=>data_re_out(1312),
            data_re_out(42)=>data_re_out(1344),
            data_re_out(43)=>data_re_out(1376),
            data_re_out(44)=>data_re_out(1408),
            data_re_out(45)=>data_re_out(1440),
            data_re_out(46)=>data_re_out(1472),
            data_re_out(47)=>data_re_out(1504),
            data_re_out(48)=>data_re_out(1536),
            data_re_out(49)=>data_re_out(1568),
            data_re_out(50)=>data_re_out(1600),
            data_re_out(51)=>data_re_out(1632),
            data_re_out(52)=>data_re_out(1664),
            data_re_out(53)=>data_re_out(1696),
            data_re_out(54)=>data_re_out(1728),
            data_re_out(55)=>data_re_out(1760),
            data_re_out(56)=>data_re_out(1792),
            data_re_out(57)=>data_re_out(1824),
            data_re_out(58)=>data_re_out(1856),
            data_re_out(59)=>data_re_out(1888),
            data_re_out(60)=>data_re_out(1920),
            data_re_out(61)=>data_re_out(1952),
            data_re_out(62)=>data_re_out(1984),
            data_re_out(63)=>data_re_out(2016),
            data_im_out(0)=>data_im_out(0),
            data_im_out(1)=>data_im_out(32),
            data_im_out(2)=>data_im_out(64),
            data_im_out(3)=>data_im_out(96),
            data_im_out(4)=>data_im_out(128),
            data_im_out(5)=>data_im_out(160),
            data_im_out(6)=>data_im_out(192),
            data_im_out(7)=>data_im_out(224),
            data_im_out(8)=>data_im_out(256),
            data_im_out(9)=>data_im_out(288),
            data_im_out(10)=>data_im_out(320),
            data_im_out(11)=>data_im_out(352),
            data_im_out(12)=>data_im_out(384),
            data_im_out(13)=>data_im_out(416),
            data_im_out(14)=>data_im_out(448),
            data_im_out(15)=>data_im_out(480),
            data_im_out(16)=>data_im_out(512),
            data_im_out(17)=>data_im_out(544),
            data_im_out(18)=>data_im_out(576),
            data_im_out(19)=>data_im_out(608),
            data_im_out(20)=>data_im_out(640),
            data_im_out(21)=>data_im_out(672),
            data_im_out(22)=>data_im_out(704),
            data_im_out(23)=>data_im_out(736),
            data_im_out(24)=>data_im_out(768),
            data_im_out(25)=>data_im_out(800),
            data_im_out(26)=>data_im_out(832),
            data_im_out(27)=>data_im_out(864),
            data_im_out(28)=>data_im_out(896),
            data_im_out(29)=>data_im_out(928),
            data_im_out(30)=>data_im_out(960),
            data_im_out(31)=>data_im_out(992),
            data_im_out(32)=>data_im_out(1024),
            data_im_out(33)=>data_im_out(1056),
            data_im_out(34)=>data_im_out(1088),
            data_im_out(35)=>data_im_out(1120),
            data_im_out(36)=>data_im_out(1152),
            data_im_out(37)=>data_im_out(1184),
            data_im_out(38)=>data_im_out(1216),
            data_im_out(39)=>data_im_out(1248),
            data_im_out(40)=>data_im_out(1280),
            data_im_out(41)=>data_im_out(1312),
            data_im_out(42)=>data_im_out(1344),
            data_im_out(43)=>data_im_out(1376),
            data_im_out(44)=>data_im_out(1408),
            data_im_out(45)=>data_im_out(1440),
            data_im_out(46)=>data_im_out(1472),
            data_im_out(47)=>data_im_out(1504),
            data_im_out(48)=>data_im_out(1536),
            data_im_out(49)=>data_im_out(1568),
            data_im_out(50)=>data_im_out(1600),
            data_im_out(51)=>data_im_out(1632),
            data_im_out(52)=>data_im_out(1664),
            data_im_out(53)=>data_im_out(1696),
            data_im_out(54)=>data_im_out(1728),
            data_im_out(55)=>data_im_out(1760),
            data_im_out(56)=>data_im_out(1792),
            data_im_out(57)=>data_im_out(1824),
            data_im_out(58)=>data_im_out(1856),
            data_im_out(59)=>data_im_out(1888),
            data_im_out(60)=>data_im_out(1920),
            data_im_out(61)=>data_im_out(1952),
            data_im_out(62)=>data_im_out(1984),
            data_im_out(63)=>data_im_out(2016)
        );           

    URFFT_PT64_1 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(1),
            data_re_in(1)=>mul_re_out(33),
            data_re_in(2)=>mul_re_out(65),
            data_re_in(3)=>mul_re_out(97),
            data_re_in(4)=>mul_re_out(129),
            data_re_in(5)=>mul_re_out(161),
            data_re_in(6)=>mul_re_out(193),
            data_re_in(7)=>mul_re_out(225),
            data_re_in(8)=>mul_re_out(257),
            data_re_in(9)=>mul_re_out(289),
            data_re_in(10)=>mul_re_out(321),
            data_re_in(11)=>mul_re_out(353),
            data_re_in(12)=>mul_re_out(385),
            data_re_in(13)=>mul_re_out(417),
            data_re_in(14)=>mul_re_out(449),
            data_re_in(15)=>mul_re_out(481),
            data_re_in(16)=>mul_re_out(513),
            data_re_in(17)=>mul_re_out(545),
            data_re_in(18)=>mul_re_out(577),
            data_re_in(19)=>mul_re_out(609),
            data_re_in(20)=>mul_re_out(641),
            data_re_in(21)=>mul_re_out(673),
            data_re_in(22)=>mul_re_out(705),
            data_re_in(23)=>mul_re_out(737),
            data_re_in(24)=>mul_re_out(769),
            data_re_in(25)=>mul_re_out(801),
            data_re_in(26)=>mul_re_out(833),
            data_re_in(27)=>mul_re_out(865),
            data_re_in(28)=>mul_re_out(897),
            data_re_in(29)=>mul_re_out(929),
            data_re_in(30)=>mul_re_out(961),
            data_re_in(31)=>mul_re_out(993),
            data_re_in(32)=>mul_re_out(1025),
            data_re_in(33)=>mul_re_out(1057),
            data_re_in(34)=>mul_re_out(1089),
            data_re_in(35)=>mul_re_out(1121),
            data_re_in(36)=>mul_re_out(1153),
            data_re_in(37)=>mul_re_out(1185),
            data_re_in(38)=>mul_re_out(1217),
            data_re_in(39)=>mul_re_out(1249),
            data_re_in(40)=>mul_re_out(1281),
            data_re_in(41)=>mul_re_out(1313),
            data_re_in(42)=>mul_re_out(1345),
            data_re_in(43)=>mul_re_out(1377),
            data_re_in(44)=>mul_re_out(1409),
            data_re_in(45)=>mul_re_out(1441),
            data_re_in(46)=>mul_re_out(1473),
            data_re_in(47)=>mul_re_out(1505),
            data_re_in(48)=>mul_re_out(1537),
            data_re_in(49)=>mul_re_out(1569),
            data_re_in(50)=>mul_re_out(1601),
            data_re_in(51)=>mul_re_out(1633),
            data_re_in(52)=>mul_re_out(1665),
            data_re_in(53)=>mul_re_out(1697),
            data_re_in(54)=>mul_re_out(1729),
            data_re_in(55)=>mul_re_out(1761),
            data_re_in(56)=>mul_re_out(1793),
            data_re_in(57)=>mul_re_out(1825),
            data_re_in(58)=>mul_re_out(1857),
            data_re_in(59)=>mul_re_out(1889),
            data_re_in(60)=>mul_re_out(1921),
            data_re_in(61)=>mul_re_out(1953),
            data_re_in(62)=>mul_re_out(1985),
            data_re_in(63)=>mul_re_out(2017),
            data_im_in(0)=>mul_im_out(1),
            data_im_in(1)=>mul_im_out(33),
            data_im_in(2)=>mul_im_out(65),
            data_im_in(3)=>mul_im_out(97),
            data_im_in(4)=>mul_im_out(129),
            data_im_in(5)=>mul_im_out(161),
            data_im_in(6)=>mul_im_out(193),
            data_im_in(7)=>mul_im_out(225),
            data_im_in(8)=>mul_im_out(257),
            data_im_in(9)=>mul_im_out(289),
            data_im_in(10)=>mul_im_out(321),
            data_im_in(11)=>mul_im_out(353),
            data_im_in(12)=>mul_im_out(385),
            data_im_in(13)=>mul_im_out(417),
            data_im_in(14)=>mul_im_out(449),
            data_im_in(15)=>mul_im_out(481),
            data_im_in(16)=>mul_im_out(513),
            data_im_in(17)=>mul_im_out(545),
            data_im_in(18)=>mul_im_out(577),
            data_im_in(19)=>mul_im_out(609),
            data_im_in(20)=>mul_im_out(641),
            data_im_in(21)=>mul_im_out(673),
            data_im_in(22)=>mul_im_out(705),
            data_im_in(23)=>mul_im_out(737),
            data_im_in(24)=>mul_im_out(769),
            data_im_in(25)=>mul_im_out(801),
            data_im_in(26)=>mul_im_out(833),
            data_im_in(27)=>mul_im_out(865),
            data_im_in(28)=>mul_im_out(897),
            data_im_in(29)=>mul_im_out(929),
            data_im_in(30)=>mul_im_out(961),
            data_im_in(31)=>mul_im_out(993),
            data_im_in(32)=>mul_im_out(1025),
            data_im_in(33)=>mul_im_out(1057),
            data_im_in(34)=>mul_im_out(1089),
            data_im_in(35)=>mul_im_out(1121),
            data_im_in(36)=>mul_im_out(1153),
            data_im_in(37)=>mul_im_out(1185),
            data_im_in(38)=>mul_im_out(1217),
            data_im_in(39)=>mul_im_out(1249),
            data_im_in(40)=>mul_im_out(1281),
            data_im_in(41)=>mul_im_out(1313),
            data_im_in(42)=>mul_im_out(1345),
            data_im_in(43)=>mul_im_out(1377),
            data_im_in(44)=>mul_im_out(1409),
            data_im_in(45)=>mul_im_out(1441),
            data_im_in(46)=>mul_im_out(1473),
            data_im_in(47)=>mul_im_out(1505),
            data_im_in(48)=>mul_im_out(1537),
            data_im_in(49)=>mul_im_out(1569),
            data_im_in(50)=>mul_im_out(1601),
            data_im_in(51)=>mul_im_out(1633),
            data_im_in(52)=>mul_im_out(1665),
            data_im_in(53)=>mul_im_out(1697),
            data_im_in(54)=>mul_im_out(1729),
            data_im_in(55)=>mul_im_out(1761),
            data_im_in(56)=>mul_im_out(1793),
            data_im_in(57)=>mul_im_out(1825),
            data_im_in(58)=>mul_im_out(1857),
            data_im_in(59)=>mul_im_out(1889),
            data_im_in(60)=>mul_im_out(1921),
            data_im_in(61)=>mul_im_out(1953),
            data_im_in(62)=>mul_im_out(1985),
            data_im_in(63)=>mul_im_out(2017),
            data_re_out(0)=>data_re_out(1),
            data_re_out(1)=>data_re_out(33),
            data_re_out(2)=>data_re_out(65),
            data_re_out(3)=>data_re_out(97),
            data_re_out(4)=>data_re_out(129),
            data_re_out(5)=>data_re_out(161),
            data_re_out(6)=>data_re_out(193),
            data_re_out(7)=>data_re_out(225),
            data_re_out(8)=>data_re_out(257),
            data_re_out(9)=>data_re_out(289),
            data_re_out(10)=>data_re_out(321),
            data_re_out(11)=>data_re_out(353),
            data_re_out(12)=>data_re_out(385),
            data_re_out(13)=>data_re_out(417),
            data_re_out(14)=>data_re_out(449),
            data_re_out(15)=>data_re_out(481),
            data_re_out(16)=>data_re_out(513),
            data_re_out(17)=>data_re_out(545),
            data_re_out(18)=>data_re_out(577),
            data_re_out(19)=>data_re_out(609),
            data_re_out(20)=>data_re_out(641),
            data_re_out(21)=>data_re_out(673),
            data_re_out(22)=>data_re_out(705),
            data_re_out(23)=>data_re_out(737),
            data_re_out(24)=>data_re_out(769),
            data_re_out(25)=>data_re_out(801),
            data_re_out(26)=>data_re_out(833),
            data_re_out(27)=>data_re_out(865),
            data_re_out(28)=>data_re_out(897),
            data_re_out(29)=>data_re_out(929),
            data_re_out(30)=>data_re_out(961),
            data_re_out(31)=>data_re_out(993),
            data_re_out(32)=>data_re_out(1025),
            data_re_out(33)=>data_re_out(1057),
            data_re_out(34)=>data_re_out(1089),
            data_re_out(35)=>data_re_out(1121),
            data_re_out(36)=>data_re_out(1153),
            data_re_out(37)=>data_re_out(1185),
            data_re_out(38)=>data_re_out(1217),
            data_re_out(39)=>data_re_out(1249),
            data_re_out(40)=>data_re_out(1281),
            data_re_out(41)=>data_re_out(1313),
            data_re_out(42)=>data_re_out(1345),
            data_re_out(43)=>data_re_out(1377),
            data_re_out(44)=>data_re_out(1409),
            data_re_out(45)=>data_re_out(1441),
            data_re_out(46)=>data_re_out(1473),
            data_re_out(47)=>data_re_out(1505),
            data_re_out(48)=>data_re_out(1537),
            data_re_out(49)=>data_re_out(1569),
            data_re_out(50)=>data_re_out(1601),
            data_re_out(51)=>data_re_out(1633),
            data_re_out(52)=>data_re_out(1665),
            data_re_out(53)=>data_re_out(1697),
            data_re_out(54)=>data_re_out(1729),
            data_re_out(55)=>data_re_out(1761),
            data_re_out(56)=>data_re_out(1793),
            data_re_out(57)=>data_re_out(1825),
            data_re_out(58)=>data_re_out(1857),
            data_re_out(59)=>data_re_out(1889),
            data_re_out(60)=>data_re_out(1921),
            data_re_out(61)=>data_re_out(1953),
            data_re_out(62)=>data_re_out(1985),
            data_re_out(63)=>data_re_out(2017),
            data_im_out(0)=>data_im_out(1),
            data_im_out(1)=>data_im_out(33),
            data_im_out(2)=>data_im_out(65),
            data_im_out(3)=>data_im_out(97),
            data_im_out(4)=>data_im_out(129),
            data_im_out(5)=>data_im_out(161),
            data_im_out(6)=>data_im_out(193),
            data_im_out(7)=>data_im_out(225),
            data_im_out(8)=>data_im_out(257),
            data_im_out(9)=>data_im_out(289),
            data_im_out(10)=>data_im_out(321),
            data_im_out(11)=>data_im_out(353),
            data_im_out(12)=>data_im_out(385),
            data_im_out(13)=>data_im_out(417),
            data_im_out(14)=>data_im_out(449),
            data_im_out(15)=>data_im_out(481),
            data_im_out(16)=>data_im_out(513),
            data_im_out(17)=>data_im_out(545),
            data_im_out(18)=>data_im_out(577),
            data_im_out(19)=>data_im_out(609),
            data_im_out(20)=>data_im_out(641),
            data_im_out(21)=>data_im_out(673),
            data_im_out(22)=>data_im_out(705),
            data_im_out(23)=>data_im_out(737),
            data_im_out(24)=>data_im_out(769),
            data_im_out(25)=>data_im_out(801),
            data_im_out(26)=>data_im_out(833),
            data_im_out(27)=>data_im_out(865),
            data_im_out(28)=>data_im_out(897),
            data_im_out(29)=>data_im_out(929),
            data_im_out(30)=>data_im_out(961),
            data_im_out(31)=>data_im_out(993),
            data_im_out(32)=>data_im_out(1025),
            data_im_out(33)=>data_im_out(1057),
            data_im_out(34)=>data_im_out(1089),
            data_im_out(35)=>data_im_out(1121),
            data_im_out(36)=>data_im_out(1153),
            data_im_out(37)=>data_im_out(1185),
            data_im_out(38)=>data_im_out(1217),
            data_im_out(39)=>data_im_out(1249),
            data_im_out(40)=>data_im_out(1281),
            data_im_out(41)=>data_im_out(1313),
            data_im_out(42)=>data_im_out(1345),
            data_im_out(43)=>data_im_out(1377),
            data_im_out(44)=>data_im_out(1409),
            data_im_out(45)=>data_im_out(1441),
            data_im_out(46)=>data_im_out(1473),
            data_im_out(47)=>data_im_out(1505),
            data_im_out(48)=>data_im_out(1537),
            data_im_out(49)=>data_im_out(1569),
            data_im_out(50)=>data_im_out(1601),
            data_im_out(51)=>data_im_out(1633),
            data_im_out(52)=>data_im_out(1665),
            data_im_out(53)=>data_im_out(1697),
            data_im_out(54)=>data_im_out(1729),
            data_im_out(55)=>data_im_out(1761),
            data_im_out(56)=>data_im_out(1793),
            data_im_out(57)=>data_im_out(1825),
            data_im_out(58)=>data_im_out(1857),
            data_im_out(59)=>data_im_out(1889),
            data_im_out(60)=>data_im_out(1921),
            data_im_out(61)=>data_im_out(1953),
            data_im_out(62)=>data_im_out(1985),
            data_im_out(63)=>data_im_out(2017)
        );           

    URFFT_PT64_2 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(2),
            data_re_in(1)=>mul_re_out(34),
            data_re_in(2)=>mul_re_out(66),
            data_re_in(3)=>mul_re_out(98),
            data_re_in(4)=>mul_re_out(130),
            data_re_in(5)=>mul_re_out(162),
            data_re_in(6)=>mul_re_out(194),
            data_re_in(7)=>mul_re_out(226),
            data_re_in(8)=>mul_re_out(258),
            data_re_in(9)=>mul_re_out(290),
            data_re_in(10)=>mul_re_out(322),
            data_re_in(11)=>mul_re_out(354),
            data_re_in(12)=>mul_re_out(386),
            data_re_in(13)=>mul_re_out(418),
            data_re_in(14)=>mul_re_out(450),
            data_re_in(15)=>mul_re_out(482),
            data_re_in(16)=>mul_re_out(514),
            data_re_in(17)=>mul_re_out(546),
            data_re_in(18)=>mul_re_out(578),
            data_re_in(19)=>mul_re_out(610),
            data_re_in(20)=>mul_re_out(642),
            data_re_in(21)=>mul_re_out(674),
            data_re_in(22)=>mul_re_out(706),
            data_re_in(23)=>mul_re_out(738),
            data_re_in(24)=>mul_re_out(770),
            data_re_in(25)=>mul_re_out(802),
            data_re_in(26)=>mul_re_out(834),
            data_re_in(27)=>mul_re_out(866),
            data_re_in(28)=>mul_re_out(898),
            data_re_in(29)=>mul_re_out(930),
            data_re_in(30)=>mul_re_out(962),
            data_re_in(31)=>mul_re_out(994),
            data_re_in(32)=>mul_re_out(1026),
            data_re_in(33)=>mul_re_out(1058),
            data_re_in(34)=>mul_re_out(1090),
            data_re_in(35)=>mul_re_out(1122),
            data_re_in(36)=>mul_re_out(1154),
            data_re_in(37)=>mul_re_out(1186),
            data_re_in(38)=>mul_re_out(1218),
            data_re_in(39)=>mul_re_out(1250),
            data_re_in(40)=>mul_re_out(1282),
            data_re_in(41)=>mul_re_out(1314),
            data_re_in(42)=>mul_re_out(1346),
            data_re_in(43)=>mul_re_out(1378),
            data_re_in(44)=>mul_re_out(1410),
            data_re_in(45)=>mul_re_out(1442),
            data_re_in(46)=>mul_re_out(1474),
            data_re_in(47)=>mul_re_out(1506),
            data_re_in(48)=>mul_re_out(1538),
            data_re_in(49)=>mul_re_out(1570),
            data_re_in(50)=>mul_re_out(1602),
            data_re_in(51)=>mul_re_out(1634),
            data_re_in(52)=>mul_re_out(1666),
            data_re_in(53)=>mul_re_out(1698),
            data_re_in(54)=>mul_re_out(1730),
            data_re_in(55)=>mul_re_out(1762),
            data_re_in(56)=>mul_re_out(1794),
            data_re_in(57)=>mul_re_out(1826),
            data_re_in(58)=>mul_re_out(1858),
            data_re_in(59)=>mul_re_out(1890),
            data_re_in(60)=>mul_re_out(1922),
            data_re_in(61)=>mul_re_out(1954),
            data_re_in(62)=>mul_re_out(1986),
            data_re_in(63)=>mul_re_out(2018),
            data_im_in(0)=>mul_im_out(2),
            data_im_in(1)=>mul_im_out(34),
            data_im_in(2)=>mul_im_out(66),
            data_im_in(3)=>mul_im_out(98),
            data_im_in(4)=>mul_im_out(130),
            data_im_in(5)=>mul_im_out(162),
            data_im_in(6)=>mul_im_out(194),
            data_im_in(7)=>mul_im_out(226),
            data_im_in(8)=>mul_im_out(258),
            data_im_in(9)=>mul_im_out(290),
            data_im_in(10)=>mul_im_out(322),
            data_im_in(11)=>mul_im_out(354),
            data_im_in(12)=>mul_im_out(386),
            data_im_in(13)=>mul_im_out(418),
            data_im_in(14)=>mul_im_out(450),
            data_im_in(15)=>mul_im_out(482),
            data_im_in(16)=>mul_im_out(514),
            data_im_in(17)=>mul_im_out(546),
            data_im_in(18)=>mul_im_out(578),
            data_im_in(19)=>mul_im_out(610),
            data_im_in(20)=>mul_im_out(642),
            data_im_in(21)=>mul_im_out(674),
            data_im_in(22)=>mul_im_out(706),
            data_im_in(23)=>mul_im_out(738),
            data_im_in(24)=>mul_im_out(770),
            data_im_in(25)=>mul_im_out(802),
            data_im_in(26)=>mul_im_out(834),
            data_im_in(27)=>mul_im_out(866),
            data_im_in(28)=>mul_im_out(898),
            data_im_in(29)=>mul_im_out(930),
            data_im_in(30)=>mul_im_out(962),
            data_im_in(31)=>mul_im_out(994),
            data_im_in(32)=>mul_im_out(1026),
            data_im_in(33)=>mul_im_out(1058),
            data_im_in(34)=>mul_im_out(1090),
            data_im_in(35)=>mul_im_out(1122),
            data_im_in(36)=>mul_im_out(1154),
            data_im_in(37)=>mul_im_out(1186),
            data_im_in(38)=>mul_im_out(1218),
            data_im_in(39)=>mul_im_out(1250),
            data_im_in(40)=>mul_im_out(1282),
            data_im_in(41)=>mul_im_out(1314),
            data_im_in(42)=>mul_im_out(1346),
            data_im_in(43)=>mul_im_out(1378),
            data_im_in(44)=>mul_im_out(1410),
            data_im_in(45)=>mul_im_out(1442),
            data_im_in(46)=>mul_im_out(1474),
            data_im_in(47)=>mul_im_out(1506),
            data_im_in(48)=>mul_im_out(1538),
            data_im_in(49)=>mul_im_out(1570),
            data_im_in(50)=>mul_im_out(1602),
            data_im_in(51)=>mul_im_out(1634),
            data_im_in(52)=>mul_im_out(1666),
            data_im_in(53)=>mul_im_out(1698),
            data_im_in(54)=>mul_im_out(1730),
            data_im_in(55)=>mul_im_out(1762),
            data_im_in(56)=>mul_im_out(1794),
            data_im_in(57)=>mul_im_out(1826),
            data_im_in(58)=>mul_im_out(1858),
            data_im_in(59)=>mul_im_out(1890),
            data_im_in(60)=>mul_im_out(1922),
            data_im_in(61)=>mul_im_out(1954),
            data_im_in(62)=>mul_im_out(1986),
            data_im_in(63)=>mul_im_out(2018),
            data_re_out(0)=>data_re_out(2),
            data_re_out(1)=>data_re_out(34),
            data_re_out(2)=>data_re_out(66),
            data_re_out(3)=>data_re_out(98),
            data_re_out(4)=>data_re_out(130),
            data_re_out(5)=>data_re_out(162),
            data_re_out(6)=>data_re_out(194),
            data_re_out(7)=>data_re_out(226),
            data_re_out(8)=>data_re_out(258),
            data_re_out(9)=>data_re_out(290),
            data_re_out(10)=>data_re_out(322),
            data_re_out(11)=>data_re_out(354),
            data_re_out(12)=>data_re_out(386),
            data_re_out(13)=>data_re_out(418),
            data_re_out(14)=>data_re_out(450),
            data_re_out(15)=>data_re_out(482),
            data_re_out(16)=>data_re_out(514),
            data_re_out(17)=>data_re_out(546),
            data_re_out(18)=>data_re_out(578),
            data_re_out(19)=>data_re_out(610),
            data_re_out(20)=>data_re_out(642),
            data_re_out(21)=>data_re_out(674),
            data_re_out(22)=>data_re_out(706),
            data_re_out(23)=>data_re_out(738),
            data_re_out(24)=>data_re_out(770),
            data_re_out(25)=>data_re_out(802),
            data_re_out(26)=>data_re_out(834),
            data_re_out(27)=>data_re_out(866),
            data_re_out(28)=>data_re_out(898),
            data_re_out(29)=>data_re_out(930),
            data_re_out(30)=>data_re_out(962),
            data_re_out(31)=>data_re_out(994),
            data_re_out(32)=>data_re_out(1026),
            data_re_out(33)=>data_re_out(1058),
            data_re_out(34)=>data_re_out(1090),
            data_re_out(35)=>data_re_out(1122),
            data_re_out(36)=>data_re_out(1154),
            data_re_out(37)=>data_re_out(1186),
            data_re_out(38)=>data_re_out(1218),
            data_re_out(39)=>data_re_out(1250),
            data_re_out(40)=>data_re_out(1282),
            data_re_out(41)=>data_re_out(1314),
            data_re_out(42)=>data_re_out(1346),
            data_re_out(43)=>data_re_out(1378),
            data_re_out(44)=>data_re_out(1410),
            data_re_out(45)=>data_re_out(1442),
            data_re_out(46)=>data_re_out(1474),
            data_re_out(47)=>data_re_out(1506),
            data_re_out(48)=>data_re_out(1538),
            data_re_out(49)=>data_re_out(1570),
            data_re_out(50)=>data_re_out(1602),
            data_re_out(51)=>data_re_out(1634),
            data_re_out(52)=>data_re_out(1666),
            data_re_out(53)=>data_re_out(1698),
            data_re_out(54)=>data_re_out(1730),
            data_re_out(55)=>data_re_out(1762),
            data_re_out(56)=>data_re_out(1794),
            data_re_out(57)=>data_re_out(1826),
            data_re_out(58)=>data_re_out(1858),
            data_re_out(59)=>data_re_out(1890),
            data_re_out(60)=>data_re_out(1922),
            data_re_out(61)=>data_re_out(1954),
            data_re_out(62)=>data_re_out(1986),
            data_re_out(63)=>data_re_out(2018),
            data_im_out(0)=>data_im_out(2),
            data_im_out(1)=>data_im_out(34),
            data_im_out(2)=>data_im_out(66),
            data_im_out(3)=>data_im_out(98),
            data_im_out(4)=>data_im_out(130),
            data_im_out(5)=>data_im_out(162),
            data_im_out(6)=>data_im_out(194),
            data_im_out(7)=>data_im_out(226),
            data_im_out(8)=>data_im_out(258),
            data_im_out(9)=>data_im_out(290),
            data_im_out(10)=>data_im_out(322),
            data_im_out(11)=>data_im_out(354),
            data_im_out(12)=>data_im_out(386),
            data_im_out(13)=>data_im_out(418),
            data_im_out(14)=>data_im_out(450),
            data_im_out(15)=>data_im_out(482),
            data_im_out(16)=>data_im_out(514),
            data_im_out(17)=>data_im_out(546),
            data_im_out(18)=>data_im_out(578),
            data_im_out(19)=>data_im_out(610),
            data_im_out(20)=>data_im_out(642),
            data_im_out(21)=>data_im_out(674),
            data_im_out(22)=>data_im_out(706),
            data_im_out(23)=>data_im_out(738),
            data_im_out(24)=>data_im_out(770),
            data_im_out(25)=>data_im_out(802),
            data_im_out(26)=>data_im_out(834),
            data_im_out(27)=>data_im_out(866),
            data_im_out(28)=>data_im_out(898),
            data_im_out(29)=>data_im_out(930),
            data_im_out(30)=>data_im_out(962),
            data_im_out(31)=>data_im_out(994),
            data_im_out(32)=>data_im_out(1026),
            data_im_out(33)=>data_im_out(1058),
            data_im_out(34)=>data_im_out(1090),
            data_im_out(35)=>data_im_out(1122),
            data_im_out(36)=>data_im_out(1154),
            data_im_out(37)=>data_im_out(1186),
            data_im_out(38)=>data_im_out(1218),
            data_im_out(39)=>data_im_out(1250),
            data_im_out(40)=>data_im_out(1282),
            data_im_out(41)=>data_im_out(1314),
            data_im_out(42)=>data_im_out(1346),
            data_im_out(43)=>data_im_out(1378),
            data_im_out(44)=>data_im_out(1410),
            data_im_out(45)=>data_im_out(1442),
            data_im_out(46)=>data_im_out(1474),
            data_im_out(47)=>data_im_out(1506),
            data_im_out(48)=>data_im_out(1538),
            data_im_out(49)=>data_im_out(1570),
            data_im_out(50)=>data_im_out(1602),
            data_im_out(51)=>data_im_out(1634),
            data_im_out(52)=>data_im_out(1666),
            data_im_out(53)=>data_im_out(1698),
            data_im_out(54)=>data_im_out(1730),
            data_im_out(55)=>data_im_out(1762),
            data_im_out(56)=>data_im_out(1794),
            data_im_out(57)=>data_im_out(1826),
            data_im_out(58)=>data_im_out(1858),
            data_im_out(59)=>data_im_out(1890),
            data_im_out(60)=>data_im_out(1922),
            data_im_out(61)=>data_im_out(1954),
            data_im_out(62)=>data_im_out(1986),
            data_im_out(63)=>data_im_out(2018)
        );           

    URFFT_PT64_3 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(3),
            data_re_in(1)=>mul_re_out(35),
            data_re_in(2)=>mul_re_out(67),
            data_re_in(3)=>mul_re_out(99),
            data_re_in(4)=>mul_re_out(131),
            data_re_in(5)=>mul_re_out(163),
            data_re_in(6)=>mul_re_out(195),
            data_re_in(7)=>mul_re_out(227),
            data_re_in(8)=>mul_re_out(259),
            data_re_in(9)=>mul_re_out(291),
            data_re_in(10)=>mul_re_out(323),
            data_re_in(11)=>mul_re_out(355),
            data_re_in(12)=>mul_re_out(387),
            data_re_in(13)=>mul_re_out(419),
            data_re_in(14)=>mul_re_out(451),
            data_re_in(15)=>mul_re_out(483),
            data_re_in(16)=>mul_re_out(515),
            data_re_in(17)=>mul_re_out(547),
            data_re_in(18)=>mul_re_out(579),
            data_re_in(19)=>mul_re_out(611),
            data_re_in(20)=>mul_re_out(643),
            data_re_in(21)=>mul_re_out(675),
            data_re_in(22)=>mul_re_out(707),
            data_re_in(23)=>mul_re_out(739),
            data_re_in(24)=>mul_re_out(771),
            data_re_in(25)=>mul_re_out(803),
            data_re_in(26)=>mul_re_out(835),
            data_re_in(27)=>mul_re_out(867),
            data_re_in(28)=>mul_re_out(899),
            data_re_in(29)=>mul_re_out(931),
            data_re_in(30)=>mul_re_out(963),
            data_re_in(31)=>mul_re_out(995),
            data_re_in(32)=>mul_re_out(1027),
            data_re_in(33)=>mul_re_out(1059),
            data_re_in(34)=>mul_re_out(1091),
            data_re_in(35)=>mul_re_out(1123),
            data_re_in(36)=>mul_re_out(1155),
            data_re_in(37)=>mul_re_out(1187),
            data_re_in(38)=>mul_re_out(1219),
            data_re_in(39)=>mul_re_out(1251),
            data_re_in(40)=>mul_re_out(1283),
            data_re_in(41)=>mul_re_out(1315),
            data_re_in(42)=>mul_re_out(1347),
            data_re_in(43)=>mul_re_out(1379),
            data_re_in(44)=>mul_re_out(1411),
            data_re_in(45)=>mul_re_out(1443),
            data_re_in(46)=>mul_re_out(1475),
            data_re_in(47)=>mul_re_out(1507),
            data_re_in(48)=>mul_re_out(1539),
            data_re_in(49)=>mul_re_out(1571),
            data_re_in(50)=>mul_re_out(1603),
            data_re_in(51)=>mul_re_out(1635),
            data_re_in(52)=>mul_re_out(1667),
            data_re_in(53)=>mul_re_out(1699),
            data_re_in(54)=>mul_re_out(1731),
            data_re_in(55)=>mul_re_out(1763),
            data_re_in(56)=>mul_re_out(1795),
            data_re_in(57)=>mul_re_out(1827),
            data_re_in(58)=>mul_re_out(1859),
            data_re_in(59)=>mul_re_out(1891),
            data_re_in(60)=>mul_re_out(1923),
            data_re_in(61)=>mul_re_out(1955),
            data_re_in(62)=>mul_re_out(1987),
            data_re_in(63)=>mul_re_out(2019),
            data_im_in(0)=>mul_im_out(3),
            data_im_in(1)=>mul_im_out(35),
            data_im_in(2)=>mul_im_out(67),
            data_im_in(3)=>mul_im_out(99),
            data_im_in(4)=>mul_im_out(131),
            data_im_in(5)=>mul_im_out(163),
            data_im_in(6)=>mul_im_out(195),
            data_im_in(7)=>mul_im_out(227),
            data_im_in(8)=>mul_im_out(259),
            data_im_in(9)=>mul_im_out(291),
            data_im_in(10)=>mul_im_out(323),
            data_im_in(11)=>mul_im_out(355),
            data_im_in(12)=>mul_im_out(387),
            data_im_in(13)=>mul_im_out(419),
            data_im_in(14)=>mul_im_out(451),
            data_im_in(15)=>mul_im_out(483),
            data_im_in(16)=>mul_im_out(515),
            data_im_in(17)=>mul_im_out(547),
            data_im_in(18)=>mul_im_out(579),
            data_im_in(19)=>mul_im_out(611),
            data_im_in(20)=>mul_im_out(643),
            data_im_in(21)=>mul_im_out(675),
            data_im_in(22)=>mul_im_out(707),
            data_im_in(23)=>mul_im_out(739),
            data_im_in(24)=>mul_im_out(771),
            data_im_in(25)=>mul_im_out(803),
            data_im_in(26)=>mul_im_out(835),
            data_im_in(27)=>mul_im_out(867),
            data_im_in(28)=>mul_im_out(899),
            data_im_in(29)=>mul_im_out(931),
            data_im_in(30)=>mul_im_out(963),
            data_im_in(31)=>mul_im_out(995),
            data_im_in(32)=>mul_im_out(1027),
            data_im_in(33)=>mul_im_out(1059),
            data_im_in(34)=>mul_im_out(1091),
            data_im_in(35)=>mul_im_out(1123),
            data_im_in(36)=>mul_im_out(1155),
            data_im_in(37)=>mul_im_out(1187),
            data_im_in(38)=>mul_im_out(1219),
            data_im_in(39)=>mul_im_out(1251),
            data_im_in(40)=>mul_im_out(1283),
            data_im_in(41)=>mul_im_out(1315),
            data_im_in(42)=>mul_im_out(1347),
            data_im_in(43)=>mul_im_out(1379),
            data_im_in(44)=>mul_im_out(1411),
            data_im_in(45)=>mul_im_out(1443),
            data_im_in(46)=>mul_im_out(1475),
            data_im_in(47)=>mul_im_out(1507),
            data_im_in(48)=>mul_im_out(1539),
            data_im_in(49)=>mul_im_out(1571),
            data_im_in(50)=>mul_im_out(1603),
            data_im_in(51)=>mul_im_out(1635),
            data_im_in(52)=>mul_im_out(1667),
            data_im_in(53)=>mul_im_out(1699),
            data_im_in(54)=>mul_im_out(1731),
            data_im_in(55)=>mul_im_out(1763),
            data_im_in(56)=>mul_im_out(1795),
            data_im_in(57)=>mul_im_out(1827),
            data_im_in(58)=>mul_im_out(1859),
            data_im_in(59)=>mul_im_out(1891),
            data_im_in(60)=>mul_im_out(1923),
            data_im_in(61)=>mul_im_out(1955),
            data_im_in(62)=>mul_im_out(1987),
            data_im_in(63)=>mul_im_out(2019),
            data_re_out(0)=>data_re_out(3),
            data_re_out(1)=>data_re_out(35),
            data_re_out(2)=>data_re_out(67),
            data_re_out(3)=>data_re_out(99),
            data_re_out(4)=>data_re_out(131),
            data_re_out(5)=>data_re_out(163),
            data_re_out(6)=>data_re_out(195),
            data_re_out(7)=>data_re_out(227),
            data_re_out(8)=>data_re_out(259),
            data_re_out(9)=>data_re_out(291),
            data_re_out(10)=>data_re_out(323),
            data_re_out(11)=>data_re_out(355),
            data_re_out(12)=>data_re_out(387),
            data_re_out(13)=>data_re_out(419),
            data_re_out(14)=>data_re_out(451),
            data_re_out(15)=>data_re_out(483),
            data_re_out(16)=>data_re_out(515),
            data_re_out(17)=>data_re_out(547),
            data_re_out(18)=>data_re_out(579),
            data_re_out(19)=>data_re_out(611),
            data_re_out(20)=>data_re_out(643),
            data_re_out(21)=>data_re_out(675),
            data_re_out(22)=>data_re_out(707),
            data_re_out(23)=>data_re_out(739),
            data_re_out(24)=>data_re_out(771),
            data_re_out(25)=>data_re_out(803),
            data_re_out(26)=>data_re_out(835),
            data_re_out(27)=>data_re_out(867),
            data_re_out(28)=>data_re_out(899),
            data_re_out(29)=>data_re_out(931),
            data_re_out(30)=>data_re_out(963),
            data_re_out(31)=>data_re_out(995),
            data_re_out(32)=>data_re_out(1027),
            data_re_out(33)=>data_re_out(1059),
            data_re_out(34)=>data_re_out(1091),
            data_re_out(35)=>data_re_out(1123),
            data_re_out(36)=>data_re_out(1155),
            data_re_out(37)=>data_re_out(1187),
            data_re_out(38)=>data_re_out(1219),
            data_re_out(39)=>data_re_out(1251),
            data_re_out(40)=>data_re_out(1283),
            data_re_out(41)=>data_re_out(1315),
            data_re_out(42)=>data_re_out(1347),
            data_re_out(43)=>data_re_out(1379),
            data_re_out(44)=>data_re_out(1411),
            data_re_out(45)=>data_re_out(1443),
            data_re_out(46)=>data_re_out(1475),
            data_re_out(47)=>data_re_out(1507),
            data_re_out(48)=>data_re_out(1539),
            data_re_out(49)=>data_re_out(1571),
            data_re_out(50)=>data_re_out(1603),
            data_re_out(51)=>data_re_out(1635),
            data_re_out(52)=>data_re_out(1667),
            data_re_out(53)=>data_re_out(1699),
            data_re_out(54)=>data_re_out(1731),
            data_re_out(55)=>data_re_out(1763),
            data_re_out(56)=>data_re_out(1795),
            data_re_out(57)=>data_re_out(1827),
            data_re_out(58)=>data_re_out(1859),
            data_re_out(59)=>data_re_out(1891),
            data_re_out(60)=>data_re_out(1923),
            data_re_out(61)=>data_re_out(1955),
            data_re_out(62)=>data_re_out(1987),
            data_re_out(63)=>data_re_out(2019),
            data_im_out(0)=>data_im_out(3),
            data_im_out(1)=>data_im_out(35),
            data_im_out(2)=>data_im_out(67),
            data_im_out(3)=>data_im_out(99),
            data_im_out(4)=>data_im_out(131),
            data_im_out(5)=>data_im_out(163),
            data_im_out(6)=>data_im_out(195),
            data_im_out(7)=>data_im_out(227),
            data_im_out(8)=>data_im_out(259),
            data_im_out(9)=>data_im_out(291),
            data_im_out(10)=>data_im_out(323),
            data_im_out(11)=>data_im_out(355),
            data_im_out(12)=>data_im_out(387),
            data_im_out(13)=>data_im_out(419),
            data_im_out(14)=>data_im_out(451),
            data_im_out(15)=>data_im_out(483),
            data_im_out(16)=>data_im_out(515),
            data_im_out(17)=>data_im_out(547),
            data_im_out(18)=>data_im_out(579),
            data_im_out(19)=>data_im_out(611),
            data_im_out(20)=>data_im_out(643),
            data_im_out(21)=>data_im_out(675),
            data_im_out(22)=>data_im_out(707),
            data_im_out(23)=>data_im_out(739),
            data_im_out(24)=>data_im_out(771),
            data_im_out(25)=>data_im_out(803),
            data_im_out(26)=>data_im_out(835),
            data_im_out(27)=>data_im_out(867),
            data_im_out(28)=>data_im_out(899),
            data_im_out(29)=>data_im_out(931),
            data_im_out(30)=>data_im_out(963),
            data_im_out(31)=>data_im_out(995),
            data_im_out(32)=>data_im_out(1027),
            data_im_out(33)=>data_im_out(1059),
            data_im_out(34)=>data_im_out(1091),
            data_im_out(35)=>data_im_out(1123),
            data_im_out(36)=>data_im_out(1155),
            data_im_out(37)=>data_im_out(1187),
            data_im_out(38)=>data_im_out(1219),
            data_im_out(39)=>data_im_out(1251),
            data_im_out(40)=>data_im_out(1283),
            data_im_out(41)=>data_im_out(1315),
            data_im_out(42)=>data_im_out(1347),
            data_im_out(43)=>data_im_out(1379),
            data_im_out(44)=>data_im_out(1411),
            data_im_out(45)=>data_im_out(1443),
            data_im_out(46)=>data_im_out(1475),
            data_im_out(47)=>data_im_out(1507),
            data_im_out(48)=>data_im_out(1539),
            data_im_out(49)=>data_im_out(1571),
            data_im_out(50)=>data_im_out(1603),
            data_im_out(51)=>data_im_out(1635),
            data_im_out(52)=>data_im_out(1667),
            data_im_out(53)=>data_im_out(1699),
            data_im_out(54)=>data_im_out(1731),
            data_im_out(55)=>data_im_out(1763),
            data_im_out(56)=>data_im_out(1795),
            data_im_out(57)=>data_im_out(1827),
            data_im_out(58)=>data_im_out(1859),
            data_im_out(59)=>data_im_out(1891),
            data_im_out(60)=>data_im_out(1923),
            data_im_out(61)=>data_im_out(1955),
            data_im_out(62)=>data_im_out(1987),
            data_im_out(63)=>data_im_out(2019)
        );           

    URFFT_PT64_4 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(4),
            data_re_in(1)=>mul_re_out(36),
            data_re_in(2)=>mul_re_out(68),
            data_re_in(3)=>mul_re_out(100),
            data_re_in(4)=>mul_re_out(132),
            data_re_in(5)=>mul_re_out(164),
            data_re_in(6)=>mul_re_out(196),
            data_re_in(7)=>mul_re_out(228),
            data_re_in(8)=>mul_re_out(260),
            data_re_in(9)=>mul_re_out(292),
            data_re_in(10)=>mul_re_out(324),
            data_re_in(11)=>mul_re_out(356),
            data_re_in(12)=>mul_re_out(388),
            data_re_in(13)=>mul_re_out(420),
            data_re_in(14)=>mul_re_out(452),
            data_re_in(15)=>mul_re_out(484),
            data_re_in(16)=>mul_re_out(516),
            data_re_in(17)=>mul_re_out(548),
            data_re_in(18)=>mul_re_out(580),
            data_re_in(19)=>mul_re_out(612),
            data_re_in(20)=>mul_re_out(644),
            data_re_in(21)=>mul_re_out(676),
            data_re_in(22)=>mul_re_out(708),
            data_re_in(23)=>mul_re_out(740),
            data_re_in(24)=>mul_re_out(772),
            data_re_in(25)=>mul_re_out(804),
            data_re_in(26)=>mul_re_out(836),
            data_re_in(27)=>mul_re_out(868),
            data_re_in(28)=>mul_re_out(900),
            data_re_in(29)=>mul_re_out(932),
            data_re_in(30)=>mul_re_out(964),
            data_re_in(31)=>mul_re_out(996),
            data_re_in(32)=>mul_re_out(1028),
            data_re_in(33)=>mul_re_out(1060),
            data_re_in(34)=>mul_re_out(1092),
            data_re_in(35)=>mul_re_out(1124),
            data_re_in(36)=>mul_re_out(1156),
            data_re_in(37)=>mul_re_out(1188),
            data_re_in(38)=>mul_re_out(1220),
            data_re_in(39)=>mul_re_out(1252),
            data_re_in(40)=>mul_re_out(1284),
            data_re_in(41)=>mul_re_out(1316),
            data_re_in(42)=>mul_re_out(1348),
            data_re_in(43)=>mul_re_out(1380),
            data_re_in(44)=>mul_re_out(1412),
            data_re_in(45)=>mul_re_out(1444),
            data_re_in(46)=>mul_re_out(1476),
            data_re_in(47)=>mul_re_out(1508),
            data_re_in(48)=>mul_re_out(1540),
            data_re_in(49)=>mul_re_out(1572),
            data_re_in(50)=>mul_re_out(1604),
            data_re_in(51)=>mul_re_out(1636),
            data_re_in(52)=>mul_re_out(1668),
            data_re_in(53)=>mul_re_out(1700),
            data_re_in(54)=>mul_re_out(1732),
            data_re_in(55)=>mul_re_out(1764),
            data_re_in(56)=>mul_re_out(1796),
            data_re_in(57)=>mul_re_out(1828),
            data_re_in(58)=>mul_re_out(1860),
            data_re_in(59)=>mul_re_out(1892),
            data_re_in(60)=>mul_re_out(1924),
            data_re_in(61)=>mul_re_out(1956),
            data_re_in(62)=>mul_re_out(1988),
            data_re_in(63)=>mul_re_out(2020),
            data_im_in(0)=>mul_im_out(4),
            data_im_in(1)=>mul_im_out(36),
            data_im_in(2)=>mul_im_out(68),
            data_im_in(3)=>mul_im_out(100),
            data_im_in(4)=>mul_im_out(132),
            data_im_in(5)=>mul_im_out(164),
            data_im_in(6)=>mul_im_out(196),
            data_im_in(7)=>mul_im_out(228),
            data_im_in(8)=>mul_im_out(260),
            data_im_in(9)=>mul_im_out(292),
            data_im_in(10)=>mul_im_out(324),
            data_im_in(11)=>mul_im_out(356),
            data_im_in(12)=>mul_im_out(388),
            data_im_in(13)=>mul_im_out(420),
            data_im_in(14)=>mul_im_out(452),
            data_im_in(15)=>mul_im_out(484),
            data_im_in(16)=>mul_im_out(516),
            data_im_in(17)=>mul_im_out(548),
            data_im_in(18)=>mul_im_out(580),
            data_im_in(19)=>mul_im_out(612),
            data_im_in(20)=>mul_im_out(644),
            data_im_in(21)=>mul_im_out(676),
            data_im_in(22)=>mul_im_out(708),
            data_im_in(23)=>mul_im_out(740),
            data_im_in(24)=>mul_im_out(772),
            data_im_in(25)=>mul_im_out(804),
            data_im_in(26)=>mul_im_out(836),
            data_im_in(27)=>mul_im_out(868),
            data_im_in(28)=>mul_im_out(900),
            data_im_in(29)=>mul_im_out(932),
            data_im_in(30)=>mul_im_out(964),
            data_im_in(31)=>mul_im_out(996),
            data_im_in(32)=>mul_im_out(1028),
            data_im_in(33)=>mul_im_out(1060),
            data_im_in(34)=>mul_im_out(1092),
            data_im_in(35)=>mul_im_out(1124),
            data_im_in(36)=>mul_im_out(1156),
            data_im_in(37)=>mul_im_out(1188),
            data_im_in(38)=>mul_im_out(1220),
            data_im_in(39)=>mul_im_out(1252),
            data_im_in(40)=>mul_im_out(1284),
            data_im_in(41)=>mul_im_out(1316),
            data_im_in(42)=>mul_im_out(1348),
            data_im_in(43)=>mul_im_out(1380),
            data_im_in(44)=>mul_im_out(1412),
            data_im_in(45)=>mul_im_out(1444),
            data_im_in(46)=>mul_im_out(1476),
            data_im_in(47)=>mul_im_out(1508),
            data_im_in(48)=>mul_im_out(1540),
            data_im_in(49)=>mul_im_out(1572),
            data_im_in(50)=>mul_im_out(1604),
            data_im_in(51)=>mul_im_out(1636),
            data_im_in(52)=>mul_im_out(1668),
            data_im_in(53)=>mul_im_out(1700),
            data_im_in(54)=>mul_im_out(1732),
            data_im_in(55)=>mul_im_out(1764),
            data_im_in(56)=>mul_im_out(1796),
            data_im_in(57)=>mul_im_out(1828),
            data_im_in(58)=>mul_im_out(1860),
            data_im_in(59)=>mul_im_out(1892),
            data_im_in(60)=>mul_im_out(1924),
            data_im_in(61)=>mul_im_out(1956),
            data_im_in(62)=>mul_im_out(1988),
            data_im_in(63)=>mul_im_out(2020),
            data_re_out(0)=>data_re_out(4),
            data_re_out(1)=>data_re_out(36),
            data_re_out(2)=>data_re_out(68),
            data_re_out(3)=>data_re_out(100),
            data_re_out(4)=>data_re_out(132),
            data_re_out(5)=>data_re_out(164),
            data_re_out(6)=>data_re_out(196),
            data_re_out(7)=>data_re_out(228),
            data_re_out(8)=>data_re_out(260),
            data_re_out(9)=>data_re_out(292),
            data_re_out(10)=>data_re_out(324),
            data_re_out(11)=>data_re_out(356),
            data_re_out(12)=>data_re_out(388),
            data_re_out(13)=>data_re_out(420),
            data_re_out(14)=>data_re_out(452),
            data_re_out(15)=>data_re_out(484),
            data_re_out(16)=>data_re_out(516),
            data_re_out(17)=>data_re_out(548),
            data_re_out(18)=>data_re_out(580),
            data_re_out(19)=>data_re_out(612),
            data_re_out(20)=>data_re_out(644),
            data_re_out(21)=>data_re_out(676),
            data_re_out(22)=>data_re_out(708),
            data_re_out(23)=>data_re_out(740),
            data_re_out(24)=>data_re_out(772),
            data_re_out(25)=>data_re_out(804),
            data_re_out(26)=>data_re_out(836),
            data_re_out(27)=>data_re_out(868),
            data_re_out(28)=>data_re_out(900),
            data_re_out(29)=>data_re_out(932),
            data_re_out(30)=>data_re_out(964),
            data_re_out(31)=>data_re_out(996),
            data_re_out(32)=>data_re_out(1028),
            data_re_out(33)=>data_re_out(1060),
            data_re_out(34)=>data_re_out(1092),
            data_re_out(35)=>data_re_out(1124),
            data_re_out(36)=>data_re_out(1156),
            data_re_out(37)=>data_re_out(1188),
            data_re_out(38)=>data_re_out(1220),
            data_re_out(39)=>data_re_out(1252),
            data_re_out(40)=>data_re_out(1284),
            data_re_out(41)=>data_re_out(1316),
            data_re_out(42)=>data_re_out(1348),
            data_re_out(43)=>data_re_out(1380),
            data_re_out(44)=>data_re_out(1412),
            data_re_out(45)=>data_re_out(1444),
            data_re_out(46)=>data_re_out(1476),
            data_re_out(47)=>data_re_out(1508),
            data_re_out(48)=>data_re_out(1540),
            data_re_out(49)=>data_re_out(1572),
            data_re_out(50)=>data_re_out(1604),
            data_re_out(51)=>data_re_out(1636),
            data_re_out(52)=>data_re_out(1668),
            data_re_out(53)=>data_re_out(1700),
            data_re_out(54)=>data_re_out(1732),
            data_re_out(55)=>data_re_out(1764),
            data_re_out(56)=>data_re_out(1796),
            data_re_out(57)=>data_re_out(1828),
            data_re_out(58)=>data_re_out(1860),
            data_re_out(59)=>data_re_out(1892),
            data_re_out(60)=>data_re_out(1924),
            data_re_out(61)=>data_re_out(1956),
            data_re_out(62)=>data_re_out(1988),
            data_re_out(63)=>data_re_out(2020),
            data_im_out(0)=>data_im_out(4),
            data_im_out(1)=>data_im_out(36),
            data_im_out(2)=>data_im_out(68),
            data_im_out(3)=>data_im_out(100),
            data_im_out(4)=>data_im_out(132),
            data_im_out(5)=>data_im_out(164),
            data_im_out(6)=>data_im_out(196),
            data_im_out(7)=>data_im_out(228),
            data_im_out(8)=>data_im_out(260),
            data_im_out(9)=>data_im_out(292),
            data_im_out(10)=>data_im_out(324),
            data_im_out(11)=>data_im_out(356),
            data_im_out(12)=>data_im_out(388),
            data_im_out(13)=>data_im_out(420),
            data_im_out(14)=>data_im_out(452),
            data_im_out(15)=>data_im_out(484),
            data_im_out(16)=>data_im_out(516),
            data_im_out(17)=>data_im_out(548),
            data_im_out(18)=>data_im_out(580),
            data_im_out(19)=>data_im_out(612),
            data_im_out(20)=>data_im_out(644),
            data_im_out(21)=>data_im_out(676),
            data_im_out(22)=>data_im_out(708),
            data_im_out(23)=>data_im_out(740),
            data_im_out(24)=>data_im_out(772),
            data_im_out(25)=>data_im_out(804),
            data_im_out(26)=>data_im_out(836),
            data_im_out(27)=>data_im_out(868),
            data_im_out(28)=>data_im_out(900),
            data_im_out(29)=>data_im_out(932),
            data_im_out(30)=>data_im_out(964),
            data_im_out(31)=>data_im_out(996),
            data_im_out(32)=>data_im_out(1028),
            data_im_out(33)=>data_im_out(1060),
            data_im_out(34)=>data_im_out(1092),
            data_im_out(35)=>data_im_out(1124),
            data_im_out(36)=>data_im_out(1156),
            data_im_out(37)=>data_im_out(1188),
            data_im_out(38)=>data_im_out(1220),
            data_im_out(39)=>data_im_out(1252),
            data_im_out(40)=>data_im_out(1284),
            data_im_out(41)=>data_im_out(1316),
            data_im_out(42)=>data_im_out(1348),
            data_im_out(43)=>data_im_out(1380),
            data_im_out(44)=>data_im_out(1412),
            data_im_out(45)=>data_im_out(1444),
            data_im_out(46)=>data_im_out(1476),
            data_im_out(47)=>data_im_out(1508),
            data_im_out(48)=>data_im_out(1540),
            data_im_out(49)=>data_im_out(1572),
            data_im_out(50)=>data_im_out(1604),
            data_im_out(51)=>data_im_out(1636),
            data_im_out(52)=>data_im_out(1668),
            data_im_out(53)=>data_im_out(1700),
            data_im_out(54)=>data_im_out(1732),
            data_im_out(55)=>data_im_out(1764),
            data_im_out(56)=>data_im_out(1796),
            data_im_out(57)=>data_im_out(1828),
            data_im_out(58)=>data_im_out(1860),
            data_im_out(59)=>data_im_out(1892),
            data_im_out(60)=>data_im_out(1924),
            data_im_out(61)=>data_im_out(1956),
            data_im_out(62)=>data_im_out(1988),
            data_im_out(63)=>data_im_out(2020)
        );           

    URFFT_PT64_5 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(5),
            data_re_in(1)=>mul_re_out(37),
            data_re_in(2)=>mul_re_out(69),
            data_re_in(3)=>mul_re_out(101),
            data_re_in(4)=>mul_re_out(133),
            data_re_in(5)=>mul_re_out(165),
            data_re_in(6)=>mul_re_out(197),
            data_re_in(7)=>mul_re_out(229),
            data_re_in(8)=>mul_re_out(261),
            data_re_in(9)=>mul_re_out(293),
            data_re_in(10)=>mul_re_out(325),
            data_re_in(11)=>mul_re_out(357),
            data_re_in(12)=>mul_re_out(389),
            data_re_in(13)=>mul_re_out(421),
            data_re_in(14)=>mul_re_out(453),
            data_re_in(15)=>mul_re_out(485),
            data_re_in(16)=>mul_re_out(517),
            data_re_in(17)=>mul_re_out(549),
            data_re_in(18)=>mul_re_out(581),
            data_re_in(19)=>mul_re_out(613),
            data_re_in(20)=>mul_re_out(645),
            data_re_in(21)=>mul_re_out(677),
            data_re_in(22)=>mul_re_out(709),
            data_re_in(23)=>mul_re_out(741),
            data_re_in(24)=>mul_re_out(773),
            data_re_in(25)=>mul_re_out(805),
            data_re_in(26)=>mul_re_out(837),
            data_re_in(27)=>mul_re_out(869),
            data_re_in(28)=>mul_re_out(901),
            data_re_in(29)=>mul_re_out(933),
            data_re_in(30)=>mul_re_out(965),
            data_re_in(31)=>mul_re_out(997),
            data_re_in(32)=>mul_re_out(1029),
            data_re_in(33)=>mul_re_out(1061),
            data_re_in(34)=>mul_re_out(1093),
            data_re_in(35)=>mul_re_out(1125),
            data_re_in(36)=>mul_re_out(1157),
            data_re_in(37)=>mul_re_out(1189),
            data_re_in(38)=>mul_re_out(1221),
            data_re_in(39)=>mul_re_out(1253),
            data_re_in(40)=>mul_re_out(1285),
            data_re_in(41)=>mul_re_out(1317),
            data_re_in(42)=>mul_re_out(1349),
            data_re_in(43)=>mul_re_out(1381),
            data_re_in(44)=>mul_re_out(1413),
            data_re_in(45)=>mul_re_out(1445),
            data_re_in(46)=>mul_re_out(1477),
            data_re_in(47)=>mul_re_out(1509),
            data_re_in(48)=>mul_re_out(1541),
            data_re_in(49)=>mul_re_out(1573),
            data_re_in(50)=>mul_re_out(1605),
            data_re_in(51)=>mul_re_out(1637),
            data_re_in(52)=>mul_re_out(1669),
            data_re_in(53)=>mul_re_out(1701),
            data_re_in(54)=>mul_re_out(1733),
            data_re_in(55)=>mul_re_out(1765),
            data_re_in(56)=>mul_re_out(1797),
            data_re_in(57)=>mul_re_out(1829),
            data_re_in(58)=>mul_re_out(1861),
            data_re_in(59)=>mul_re_out(1893),
            data_re_in(60)=>mul_re_out(1925),
            data_re_in(61)=>mul_re_out(1957),
            data_re_in(62)=>mul_re_out(1989),
            data_re_in(63)=>mul_re_out(2021),
            data_im_in(0)=>mul_im_out(5),
            data_im_in(1)=>mul_im_out(37),
            data_im_in(2)=>mul_im_out(69),
            data_im_in(3)=>mul_im_out(101),
            data_im_in(4)=>mul_im_out(133),
            data_im_in(5)=>mul_im_out(165),
            data_im_in(6)=>mul_im_out(197),
            data_im_in(7)=>mul_im_out(229),
            data_im_in(8)=>mul_im_out(261),
            data_im_in(9)=>mul_im_out(293),
            data_im_in(10)=>mul_im_out(325),
            data_im_in(11)=>mul_im_out(357),
            data_im_in(12)=>mul_im_out(389),
            data_im_in(13)=>mul_im_out(421),
            data_im_in(14)=>mul_im_out(453),
            data_im_in(15)=>mul_im_out(485),
            data_im_in(16)=>mul_im_out(517),
            data_im_in(17)=>mul_im_out(549),
            data_im_in(18)=>mul_im_out(581),
            data_im_in(19)=>mul_im_out(613),
            data_im_in(20)=>mul_im_out(645),
            data_im_in(21)=>mul_im_out(677),
            data_im_in(22)=>mul_im_out(709),
            data_im_in(23)=>mul_im_out(741),
            data_im_in(24)=>mul_im_out(773),
            data_im_in(25)=>mul_im_out(805),
            data_im_in(26)=>mul_im_out(837),
            data_im_in(27)=>mul_im_out(869),
            data_im_in(28)=>mul_im_out(901),
            data_im_in(29)=>mul_im_out(933),
            data_im_in(30)=>mul_im_out(965),
            data_im_in(31)=>mul_im_out(997),
            data_im_in(32)=>mul_im_out(1029),
            data_im_in(33)=>mul_im_out(1061),
            data_im_in(34)=>mul_im_out(1093),
            data_im_in(35)=>mul_im_out(1125),
            data_im_in(36)=>mul_im_out(1157),
            data_im_in(37)=>mul_im_out(1189),
            data_im_in(38)=>mul_im_out(1221),
            data_im_in(39)=>mul_im_out(1253),
            data_im_in(40)=>mul_im_out(1285),
            data_im_in(41)=>mul_im_out(1317),
            data_im_in(42)=>mul_im_out(1349),
            data_im_in(43)=>mul_im_out(1381),
            data_im_in(44)=>mul_im_out(1413),
            data_im_in(45)=>mul_im_out(1445),
            data_im_in(46)=>mul_im_out(1477),
            data_im_in(47)=>mul_im_out(1509),
            data_im_in(48)=>mul_im_out(1541),
            data_im_in(49)=>mul_im_out(1573),
            data_im_in(50)=>mul_im_out(1605),
            data_im_in(51)=>mul_im_out(1637),
            data_im_in(52)=>mul_im_out(1669),
            data_im_in(53)=>mul_im_out(1701),
            data_im_in(54)=>mul_im_out(1733),
            data_im_in(55)=>mul_im_out(1765),
            data_im_in(56)=>mul_im_out(1797),
            data_im_in(57)=>mul_im_out(1829),
            data_im_in(58)=>mul_im_out(1861),
            data_im_in(59)=>mul_im_out(1893),
            data_im_in(60)=>mul_im_out(1925),
            data_im_in(61)=>mul_im_out(1957),
            data_im_in(62)=>mul_im_out(1989),
            data_im_in(63)=>mul_im_out(2021),
            data_re_out(0)=>data_re_out(5),
            data_re_out(1)=>data_re_out(37),
            data_re_out(2)=>data_re_out(69),
            data_re_out(3)=>data_re_out(101),
            data_re_out(4)=>data_re_out(133),
            data_re_out(5)=>data_re_out(165),
            data_re_out(6)=>data_re_out(197),
            data_re_out(7)=>data_re_out(229),
            data_re_out(8)=>data_re_out(261),
            data_re_out(9)=>data_re_out(293),
            data_re_out(10)=>data_re_out(325),
            data_re_out(11)=>data_re_out(357),
            data_re_out(12)=>data_re_out(389),
            data_re_out(13)=>data_re_out(421),
            data_re_out(14)=>data_re_out(453),
            data_re_out(15)=>data_re_out(485),
            data_re_out(16)=>data_re_out(517),
            data_re_out(17)=>data_re_out(549),
            data_re_out(18)=>data_re_out(581),
            data_re_out(19)=>data_re_out(613),
            data_re_out(20)=>data_re_out(645),
            data_re_out(21)=>data_re_out(677),
            data_re_out(22)=>data_re_out(709),
            data_re_out(23)=>data_re_out(741),
            data_re_out(24)=>data_re_out(773),
            data_re_out(25)=>data_re_out(805),
            data_re_out(26)=>data_re_out(837),
            data_re_out(27)=>data_re_out(869),
            data_re_out(28)=>data_re_out(901),
            data_re_out(29)=>data_re_out(933),
            data_re_out(30)=>data_re_out(965),
            data_re_out(31)=>data_re_out(997),
            data_re_out(32)=>data_re_out(1029),
            data_re_out(33)=>data_re_out(1061),
            data_re_out(34)=>data_re_out(1093),
            data_re_out(35)=>data_re_out(1125),
            data_re_out(36)=>data_re_out(1157),
            data_re_out(37)=>data_re_out(1189),
            data_re_out(38)=>data_re_out(1221),
            data_re_out(39)=>data_re_out(1253),
            data_re_out(40)=>data_re_out(1285),
            data_re_out(41)=>data_re_out(1317),
            data_re_out(42)=>data_re_out(1349),
            data_re_out(43)=>data_re_out(1381),
            data_re_out(44)=>data_re_out(1413),
            data_re_out(45)=>data_re_out(1445),
            data_re_out(46)=>data_re_out(1477),
            data_re_out(47)=>data_re_out(1509),
            data_re_out(48)=>data_re_out(1541),
            data_re_out(49)=>data_re_out(1573),
            data_re_out(50)=>data_re_out(1605),
            data_re_out(51)=>data_re_out(1637),
            data_re_out(52)=>data_re_out(1669),
            data_re_out(53)=>data_re_out(1701),
            data_re_out(54)=>data_re_out(1733),
            data_re_out(55)=>data_re_out(1765),
            data_re_out(56)=>data_re_out(1797),
            data_re_out(57)=>data_re_out(1829),
            data_re_out(58)=>data_re_out(1861),
            data_re_out(59)=>data_re_out(1893),
            data_re_out(60)=>data_re_out(1925),
            data_re_out(61)=>data_re_out(1957),
            data_re_out(62)=>data_re_out(1989),
            data_re_out(63)=>data_re_out(2021),
            data_im_out(0)=>data_im_out(5),
            data_im_out(1)=>data_im_out(37),
            data_im_out(2)=>data_im_out(69),
            data_im_out(3)=>data_im_out(101),
            data_im_out(4)=>data_im_out(133),
            data_im_out(5)=>data_im_out(165),
            data_im_out(6)=>data_im_out(197),
            data_im_out(7)=>data_im_out(229),
            data_im_out(8)=>data_im_out(261),
            data_im_out(9)=>data_im_out(293),
            data_im_out(10)=>data_im_out(325),
            data_im_out(11)=>data_im_out(357),
            data_im_out(12)=>data_im_out(389),
            data_im_out(13)=>data_im_out(421),
            data_im_out(14)=>data_im_out(453),
            data_im_out(15)=>data_im_out(485),
            data_im_out(16)=>data_im_out(517),
            data_im_out(17)=>data_im_out(549),
            data_im_out(18)=>data_im_out(581),
            data_im_out(19)=>data_im_out(613),
            data_im_out(20)=>data_im_out(645),
            data_im_out(21)=>data_im_out(677),
            data_im_out(22)=>data_im_out(709),
            data_im_out(23)=>data_im_out(741),
            data_im_out(24)=>data_im_out(773),
            data_im_out(25)=>data_im_out(805),
            data_im_out(26)=>data_im_out(837),
            data_im_out(27)=>data_im_out(869),
            data_im_out(28)=>data_im_out(901),
            data_im_out(29)=>data_im_out(933),
            data_im_out(30)=>data_im_out(965),
            data_im_out(31)=>data_im_out(997),
            data_im_out(32)=>data_im_out(1029),
            data_im_out(33)=>data_im_out(1061),
            data_im_out(34)=>data_im_out(1093),
            data_im_out(35)=>data_im_out(1125),
            data_im_out(36)=>data_im_out(1157),
            data_im_out(37)=>data_im_out(1189),
            data_im_out(38)=>data_im_out(1221),
            data_im_out(39)=>data_im_out(1253),
            data_im_out(40)=>data_im_out(1285),
            data_im_out(41)=>data_im_out(1317),
            data_im_out(42)=>data_im_out(1349),
            data_im_out(43)=>data_im_out(1381),
            data_im_out(44)=>data_im_out(1413),
            data_im_out(45)=>data_im_out(1445),
            data_im_out(46)=>data_im_out(1477),
            data_im_out(47)=>data_im_out(1509),
            data_im_out(48)=>data_im_out(1541),
            data_im_out(49)=>data_im_out(1573),
            data_im_out(50)=>data_im_out(1605),
            data_im_out(51)=>data_im_out(1637),
            data_im_out(52)=>data_im_out(1669),
            data_im_out(53)=>data_im_out(1701),
            data_im_out(54)=>data_im_out(1733),
            data_im_out(55)=>data_im_out(1765),
            data_im_out(56)=>data_im_out(1797),
            data_im_out(57)=>data_im_out(1829),
            data_im_out(58)=>data_im_out(1861),
            data_im_out(59)=>data_im_out(1893),
            data_im_out(60)=>data_im_out(1925),
            data_im_out(61)=>data_im_out(1957),
            data_im_out(62)=>data_im_out(1989),
            data_im_out(63)=>data_im_out(2021)
        );           

    URFFT_PT64_6 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(6),
            data_re_in(1)=>mul_re_out(38),
            data_re_in(2)=>mul_re_out(70),
            data_re_in(3)=>mul_re_out(102),
            data_re_in(4)=>mul_re_out(134),
            data_re_in(5)=>mul_re_out(166),
            data_re_in(6)=>mul_re_out(198),
            data_re_in(7)=>mul_re_out(230),
            data_re_in(8)=>mul_re_out(262),
            data_re_in(9)=>mul_re_out(294),
            data_re_in(10)=>mul_re_out(326),
            data_re_in(11)=>mul_re_out(358),
            data_re_in(12)=>mul_re_out(390),
            data_re_in(13)=>mul_re_out(422),
            data_re_in(14)=>mul_re_out(454),
            data_re_in(15)=>mul_re_out(486),
            data_re_in(16)=>mul_re_out(518),
            data_re_in(17)=>mul_re_out(550),
            data_re_in(18)=>mul_re_out(582),
            data_re_in(19)=>mul_re_out(614),
            data_re_in(20)=>mul_re_out(646),
            data_re_in(21)=>mul_re_out(678),
            data_re_in(22)=>mul_re_out(710),
            data_re_in(23)=>mul_re_out(742),
            data_re_in(24)=>mul_re_out(774),
            data_re_in(25)=>mul_re_out(806),
            data_re_in(26)=>mul_re_out(838),
            data_re_in(27)=>mul_re_out(870),
            data_re_in(28)=>mul_re_out(902),
            data_re_in(29)=>mul_re_out(934),
            data_re_in(30)=>mul_re_out(966),
            data_re_in(31)=>mul_re_out(998),
            data_re_in(32)=>mul_re_out(1030),
            data_re_in(33)=>mul_re_out(1062),
            data_re_in(34)=>mul_re_out(1094),
            data_re_in(35)=>mul_re_out(1126),
            data_re_in(36)=>mul_re_out(1158),
            data_re_in(37)=>mul_re_out(1190),
            data_re_in(38)=>mul_re_out(1222),
            data_re_in(39)=>mul_re_out(1254),
            data_re_in(40)=>mul_re_out(1286),
            data_re_in(41)=>mul_re_out(1318),
            data_re_in(42)=>mul_re_out(1350),
            data_re_in(43)=>mul_re_out(1382),
            data_re_in(44)=>mul_re_out(1414),
            data_re_in(45)=>mul_re_out(1446),
            data_re_in(46)=>mul_re_out(1478),
            data_re_in(47)=>mul_re_out(1510),
            data_re_in(48)=>mul_re_out(1542),
            data_re_in(49)=>mul_re_out(1574),
            data_re_in(50)=>mul_re_out(1606),
            data_re_in(51)=>mul_re_out(1638),
            data_re_in(52)=>mul_re_out(1670),
            data_re_in(53)=>mul_re_out(1702),
            data_re_in(54)=>mul_re_out(1734),
            data_re_in(55)=>mul_re_out(1766),
            data_re_in(56)=>mul_re_out(1798),
            data_re_in(57)=>mul_re_out(1830),
            data_re_in(58)=>mul_re_out(1862),
            data_re_in(59)=>mul_re_out(1894),
            data_re_in(60)=>mul_re_out(1926),
            data_re_in(61)=>mul_re_out(1958),
            data_re_in(62)=>mul_re_out(1990),
            data_re_in(63)=>mul_re_out(2022),
            data_im_in(0)=>mul_im_out(6),
            data_im_in(1)=>mul_im_out(38),
            data_im_in(2)=>mul_im_out(70),
            data_im_in(3)=>mul_im_out(102),
            data_im_in(4)=>mul_im_out(134),
            data_im_in(5)=>mul_im_out(166),
            data_im_in(6)=>mul_im_out(198),
            data_im_in(7)=>mul_im_out(230),
            data_im_in(8)=>mul_im_out(262),
            data_im_in(9)=>mul_im_out(294),
            data_im_in(10)=>mul_im_out(326),
            data_im_in(11)=>mul_im_out(358),
            data_im_in(12)=>mul_im_out(390),
            data_im_in(13)=>mul_im_out(422),
            data_im_in(14)=>mul_im_out(454),
            data_im_in(15)=>mul_im_out(486),
            data_im_in(16)=>mul_im_out(518),
            data_im_in(17)=>mul_im_out(550),
            data_im_in(18)=>mul_im_out(582),
            data_im_in(19)=>mul_im_out(614),
            data_im_in(20)=>mul_im_out(646),
            data_im_in(21)=>mul_im_out(678),
            data_im_in(22)=>mul_im_out(710),
            data_im_in(23)=>mul_im_out(742),
            data_im_in(24)=>mul_im_out(774),
            data_im_in(25)=>mul_im_out(806),
            data_im_in(26)=>mul_im_out(838),
            data_im_in(27)=>mul_im_out(870),
            data_im_in(28)=>mul_im_out(902),
            data_im_in(29)=>mul_im_out(934),
            data_im_in(30)=>mul_im_out(966),
            data_im_in(31)=>mul_im_out(998),
            data_im_in(32)=>mul_im_out(1030),
            data_im_in(33)=>mul_im_out(1062),
            data_im_in(34)=>mul_im_out(1094),
            data_im_in(35)=>mul_im_out(1126),
            data_im_in(36)=>mul_im_out(1158),
            data_im_in(37)=>mul_im_out(1190),
            data_im_in(38)=>mul_im_out(1222),
            data_im_in(39)=>mul_im_out(1254),
            data_im_in(40)=>mul_im_out(1286),
            data_im_in(41)=>mul_im_out(1318),
            data_im_in(42)=>mul_im_out(1350),
            data_im_in(43)=>mul_im_out(1382),
            data_im_in(44)=>mul_im_out(1414),
            data_im_in(45)=>mul_im_out(1446),
            data_im_in(46)=>mul_im_out(1478),
            data_im_in(47)=>mul_im_out(1510),
            data_im_in(48)=>mul_im_out(1542),
            data_im_in(49)=>mul_im_out(1574),
            data_im_in(50)=>mul_im_out(1606),
            data_im_in(51)=>mul_im_out(1638),
            data_im_in(52)=>mul_im_out(1670),
            data_im_in(53)=>mul_im_out(1702),
            data_im_in(54)=>mul_im_out(1734),
            data_im_in(55)=>mul_im_out(1766),
            data_im_in(56)=>mul_im_out(1798),
            data_im_in(57)=>mul_im_out(1830),
            data_im_in(58)=>mul_im_out(1862),
            data_im_in(59)=>mul_im_out(1894),
            data_im_in(60)=>mul_im_out(1926),
            data_im_in(61)=>mul_im_out(1958),
            data_im_in(62)=>mul_im_out(1990),
            data_im_in(63)=>mul_im_out(2022),
            data_re_out(0)=>data_re_out(6),
            data_re_out(1)=>data_re_out(38),
            data_re_out(2)=>data_re_out(70),
            data_re_out(3)=>data_re_out(102),
            data_re_out(4)=>data_re_out(134),
            data_re_out(5)=>data_re_out(166),
            data_re_out(6)=>data_re_out(198),
            data_re_out(7)=>data_re_out(230),
            data_re_out(8)=>data_re_out(262),
            data_re_out(9)=>data_re_out(294),
            data_re_out(10)=>data_re_out(326),
            data_re_out(11)=>data_re_out(358),
            data_re_out(12)=>data_re_out(390),
            data_re_out(13)=>data_re_out(422),
            data_re_out(14)=>data_re_out(454),
            data_re_out(15)=>data_re_out(486),
            data_re_out(16)=>data_re_out(518),
            data_re_out(17)=>data_re_out(550),
            data_re_out(18)=>data_re_out(582),
            data_re_out(19)=>data_re_out(614),
            data_re_out(20)=>data_re_out(646),
            data_re_out(21)=>data_re_out(678),
            data_re_out(22)=>data_re_out(710),
            data_re_out(23)=>data_re_out(742),
            data_re_out(24)=>data_re_out(774),
            data_re_out(25)=>data_re_out(806),
            data_re_out(26)=>data_re_out(838),
            data_re_out(27)=>data_re_out(870),
            data_re_out(28)=>data_re_out(902),
            data_re_out(29)=>data_re_out(934),
            data_re_out(30)=>data_re_out(966),
            data_re_out(31)=>data_re_out(998),
            data_re_out(32)=>data_re_out(1030),
            data_re_out(33)=>data_re_out(1062),
            data_re_out(34)=>data_re_out(1094),
            data_re_out(35)=>data_re_out(1126),
            data_re_out(36)=>data_re_out(1158),
            data_re_out(37)=>data_re_out(1190),
            data_re_out(38)=>data_re_out(1222),
            data_re_out(39)=>data_re_out(1254),
            data_re_out(40)=>data_re_out(1286),
            data_re_out(41)=>data_re_out(1318),
            data_re_out(42)=>data_re_out(1350),
            data_re_out(43)=>data_re_out(1382),
            data_re_out(44)=>data_re_out(1414),
            data_re_out(45)=>data_re_out(1446),
            data_re_out(46)=>data_re_out(1478),
            data_re_out(47)=>data_re_out(1510),
            data_re_out(48)=>data_re_out(1542),
            data_re_out(49)=>data_re_out(1574),
            data_re_out(50)=>data_re_out(1606),
            data_re_out(51)=>data_re_out(1638),
            data_re_out(52)=>data_re_out(1670),
            data_re_out(53)=>data_re_out(1702),
            data_re_out(54)=>data_re_out(1734),
            data_re_out(55)=>data_re_out(1766),
            data_re_out(56)=>data_re_out(1798),
            data_re_out(57)=>data_re_out(1830),
            data_re_out(58)=>data_re_out(1862),
            data_re_out(59)=>data_re_out(1894),
            data_re_out(60)=>data_re_out(1926),
            data_re_out(61)=>data_re_out(1958),
            data_re_out(62)=>data_re_out(1990),
            data_re_out(63)=>data_re_out(2022),
            data_im_out(0)=>data_im_out(6),
            data_im_out(1)=>data_im_out(38),
            data_im_out(2)=>data_im_out(70),
            data_im_out(3)=>data_im_out(102),
            data_im_out(4)=>data_im_out(134),
            data_im_out(5)=>data_im_out(166),
            data_im_out(6)=>data_im_out(198),
            data_im_out(7)=>data_im_out(230),
            data_im_out(8)=>data_im_out(262),
            data_im_out(9)=>data_im_out(294),
            data_im_out(10)=>data_im_out(326),
            data_im_out(11)=>data_im_out(358),
            data_im_out(12)=>data_im_out(390),
            data_im_out(13)=>data_im_out(422),
            data_im_out(14)=>data_im_out(454),
            data_im_out(15)=>data_im_out(486),
            data_im_out(16)=>data_im_out(518),
            data_im_out(17)=>data_im_out(550),
            data_im_out(18)=>data_im_out(582),
            data_im_out(19)=>data_im_out(614),
            data_im_out(20)=>data_im_out(646),
            data_im_out(21)=>data_im_out(678),
            data_im_out(22)=>data_im_out(710),
            data_im_out(23)=>data_im_out(742),
            data_im_out(24)=>data_im_out(774),
            data_im_out(25)=>data_im_out(806),
            data_im_out(26)=>data_im_out(838),
            data_im_out(27)=>data_im_out(870),
            data_im_out(28)=>data_im_out(902),
            data_im_out(29)=>data_im_out(934),
            data_im_out(30)=>data_im_out(966),
            data_im_out(31)=>data_im_out(998),
            data_im_out(32)=>data_im_out(1030),
            data_im_out(33)=>data_im_out(1062),
            data_im_out(34)=>data_im_out(1094),
            data_im_out(35)=>data_im_out(1126),
            data_im_out(36)=>data_im_out(1158),
            data_im_out(37)=>data_im_out(1190),
            data_im_out(38)=>data_im_out(1222),
            data_im_out(39)=>data_im_out(1254),
            data_im_out(40)=>data_im_out(1286),
            data_im_out(41)=>data_im_out(1318),
            data_im_out(42)=>data_im_out(1350),
            data_im_out(43)=>data_im_out(1382),
            data_im_out(44)=>data_im_out(1414),
            data_im_out(45)=>data_im_out(1446),
            data_im_out(46)=>data_im_out(1478),
            data_im_out(47)=>data_im_out(1510),
            data_im_out(48)=>data_im_out(1542),
            data_im_out(49)=>data_im_out(1574),
            data_im_out(50)=>data_im_out(1606),
            data_im_out(51)=>data_im_out(1638),
            data_im_out(52)=>data_im_out(1670),
            data_im_out(53)=>data_im_out(1702),
            data_im_out(54)=>data_im_out(1734),
            data_im_out(55)=>data_im_out(1766),
            data_im_out(56)=>data_im_out(1798),
            data_im_out(57)=>data_im_out(1830),
            data_im_out(58)=>data_im_out(1862),
            data_im_out(59)=>data_im_out(1894),
            data_im_out(60)=>data_im_out(1926),
            data_im_out(61)=>data_im_out(1958),
            data_im_out(62)=>data_im_out(1990),
            data_im_out(63)=>data_im_out(2022)
        );           

    URFFT_PT64_7 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(7),
            data_re_in(1)=>mul_re_out(39),
            data_re_in(2)=>mul_re_out(71),
            data_re_in(3)=>mul_re_out(103),
            data_re_in(4)=>mul_re_out(135),
            data_re_in(5)=>mul_re_out(167),
            data_re_in(6)=>mul_re_out(199),
            data_re_in(7)=>mul_re_out(231),
            data_re_in(8)=>mul_re_out(263),
            data_re_in(9)=>mul_re_out(295),
            data_re_in(10)=>mul_re_out(327),
            data_re_in(11)=>mul_re_out(359),
            data_re_in(12)=>mul_re_out(391),
            data_re_in(13)=>mul_re_out(423),
            data_re_in(14)=>mul_re_out(455),
            data_re_in(15)=>mul_re_out(487),
            data_re_in(16)=>mul_re_out(519),
            data_re_in(17)=>mul_re_out(551),
            data_re_in(18)=>mul_re_out(583),
            data_re_in(19)=>mul_re_out(615),
            data_re_in(20)=>mul_re_out(647),
            data_re_in(21)=>mul_re_out(679),
            data_re_in(22)=>mul_re_out(711),
            data_re_in(23)=>mul_re_out(743),
            data_re_in(24)=>mul_re_out(775),
            data_re_in(25)=>mul_re_out(807),
            data_re_in(26)=>mul_re_out(839),
            data_re_in(27)=>mul_re_out(871),
            data_re_in(28)=>mul_re_out(903),
            data_re_in(29)=>mul_re_out(935),
            data_re_in(30)=>mul_re_out(967),
            data_re_in(31)=>mul_re_out(999),
            data_re_in(32)=>mul_re_out(1031),
            data_re_in(33)=>mul_re_out(1063),
            data_re_in(34)=>mul_re_out(1095),
            data_re_in(35)=>mul_re_out(1127),
            data_re_in(36)=>mul_re_out(1159),
            data_re_in(37)=>mul_re_out(1191),
            data_re_in(38)=>mul_re_out(1223),
            data_re_in(39)=>mul_re_out(1255),
            data_re_in(40)=>mul_re_out(1287),
            data_re_in(41)=>mul_re_out(1319),
            data_re_in(42)=>mul_re_out(1351),
            data_re_in(43)=>mul_re_out(1383),
            data_re_in(44)=>mul_re_out(1415),
            data_re_in(45)=>mul_re_out(1447),
            data_re_in(46)=>mul_re_out(1479),
            data_re_in(47)=>mul_re_out(1511),
            data_re_in(48)=>mul_re_out(1543),
            data_re_in(49)=>mul_re_out(1575),
            data_re_in(50)=>mul_re_out(1607),
            data_re_in(51)=>mul_re_out(1639),
            data_re_in(52)=>mul_re_out(1671),
            data_re_in(53)=>mul_re_out(1703),
            data_re_in(54)=>mul_re_out(1735),
            data_re_in(55)=>mul_re_out(1767),
            data_re_in(56)=>mul_re_out(1799),
            data_re_in(57)=>mul_re_out(1831),
            data_re_in(58)=>mul_re_out(1863),
            data_re_in(59)=>mul_re_out(1895),
            data_re_in(60)=>mul_re_out(1927),
            data_re_in(61)=>mul_re_out(1959),
            data_re_in(62)=>mul_re_out(1991),
            data_re_in(63)=>mul_re_out(2023),
            data_im_in(0)=>mul_im_out(7),
            data_im_in(1)=>mul_im_out(39),
            data_im_in(2)=>mul_im_out(71),
            data_im_in(3)=>mul_im_out(103),
            data_im_in(4)=>mul_im_out(135),
            data_im_in(5)=>mul_im_out(167),
            data_im_in(6)=>mul_im_out(199),
            data_im_in(7)=>mul_im_out(231),
            data_im_in(8)=>mul_im_out(263),
            data_im_in(9)=>mul_im_out(295),
            data_im_in(10)=>mul_im_out(327),
            data_im_in(11)=>mul_im_out(359),
            data_im_in(12)=>mul_im_out(391),
            data_im_in(13)=>mul_im_out(423),
            data_im_in(14)=>mul_im_out(455),
            data_im_in(15)=>mul_im_out(487),
            data_im_in(16)=>mul_im_out(519),
            data_im_in(17)=>mul_im_out(551),
            data_im_in(18)=>mul_im_out(583),
            data_im_in(19)=>mul_im_out(615),
            data_im_in(20)=>mul_im_out(647),
            data_im_in(21)=>mul_im_out(679),
            data_im_in(22)=>mul_im_out(711),
            data_im_in(23)=>mul_im_out(743),
            data_im_in(24)=>mul_im_out(775),
            data_im_in(25)=>mul_im_out(807),
            data_im_in(26)=>mul_im_out(839),
            data_im_in(27)=>mul_im_out(871),
            data_im_in(28)=>mul_im_out(903),
            data_im_in(29)=>mul_im_out(935),
            data_im_in(30)=>mul_im_out(967),
            data_im_in(31)=>mul_im_out(999),
            data_im_in(32)=>mul_im_out(1031),
            data_im_in(33)=>mul_im_out(1063),
            data_im_in(34)=>mul_im_out(1095),
            data_im_in(35)=>mul_im_out(1127),
            data_im_in(36)=>mul_im_out(1159),
            data_im_in(37)=>mul_im_out(1191),
            data_im_in(38)=>mul_im_out(1223),
            data_im_in(39)=>mul_im_out(1255),
            data_im_in(40)=>mul_im_out(1287),
            data_im_in(41)=>mul_im_out(1319),
            data_im_in(42)=>mul_im_out(1351),
            data_im_in(43)=>mul_im_out(1383),
            data_im_in(44)=>mul_im_out(1415),
            data_im_in(45)=>mul_im_out(1447),
            data_im_in(46)=>mul_im_out(1479),
            data_im_in(47)=>mul_im_out(1511),
            data_im_in(48)=>mul_im_out(1543),
            data_im_in(49)=>mul_im_out(1575),
            data_im_in(50)=>mul_im_out(1607),
            data_im_in(51)=>mul_im_out(1639),
            data_im_in(52)=>mul_im_out(1671),
            data_im_in(53)=>mul_im_out(1703),
            data_im_in(54)=>mul_im_out(1735),
            data_im_in(55)=>mul_im_out(1767),
            data_im_in(56)=>mul_im_out(1799),
            data_im_in(57)=>mul_im_out(1831),
            data_im_in(58)=>mul_im_out(1863),
            data_im_in(59)=>mul_im_out(1895),
            data_im_in(60)=>mul_im_out(1927),
            data_im_in(61)=>mul_im_out(1959),
            data_im_in(62)=>mul_im_out(1991),
            data_im_in(63)=>mul_im_out(2023),
            data_re_out(0)=>data_re_out(7),
            data_re_out(1)=>data_re_out(39),
            data_re_out(2)=>data_re_out(71),
            data_re_out(3)=>data_re_out(103),
            data_re_out(4)=>data_re_out(135),
            data_re_out(5)=>data_re_out(167),
            data_re_out(6)=>data_re_out(199),
            data_re_out(7)=>data_re_out(231),
            data_re_out(8)=>data_re_out(263),
            data_re_out(9)=>data_re_out(295),
            data_re_out(10)=>data_re_out(327),
            data_re_out(11)=>data_re_out(359),
            data_re_out(12)=>data_re_out(391),
            data_re_out(13)=>data_re_out(423),
            data_re_out(14)=>data_re_out(455),
            data_re_out(15)=>data_re_out(487),
            data_re_out(16)=>data_re_out(519),
            data_re_out(17)=>data_re_out(551),
            data_re_out(18)=>data_re_out(583),
            data_re_out(19)=>data_re_out(615),
            data_re_out(20)=>data_re_out(647),
            data_re_out(21)=>data_re_out(679),
            data_re_out(22)=>data_re_out(711),
            data_re_out(23)=>data_re_out(743),
            data_re_out(24)=>data_re_out(775),
            data_re_out(25)=>data_re_out(807),
            data_re_out(26)=>data_re_out(839),
            data_re_out(27)=>data_re_out(871),
            data_re_out(28)=>data_re_out(903),
            data_re_out(29)=>data_re_out(935),
            data_re_out(30)=>data_re_out(967),
            data_re_out(31)=>data_re_out(999),
            data_re_out(32)=>data_re_out(1031),
            data_re_out(33)=>data_re_out(1063),
            data_re_out(34)=>data_re_out(1095),
            data_re_out(35)=>data_re_out(1127),
            data_re_out(36)=>data_re_out(1159),
            data_re_out(37)=>data_re_out(1191),
            data_re_out(38)=>data_re_out(1223),
            data_re_out(39)=>data_re_out(1255),
            data_re_out(40)=>data_re_out(1287),
            data_re_out(41)=>data_re_out(1319),
            data_re_out(42)=>data_re_out(1351),
            data_re_out(43)=>data_re_out(1383),
            data_re_out(44)=>data_re_out(1415),
            data_re_out(45)=>data_re_out(1447),
            data_re_out(46)=>data_re_out(1479),
            data_re_out(47)=>data_re_out(1511),
            data_re_out(48)=>data_re_out(1543),
            data_re_out(49)=>data_re_out(1575),
            data_re_out(50)=>data_re_out(1607),
            data_re_out(51)=>data_re_out(1639),
            data_re_out(52)=>data_re_out(1671),
            data_re_out(53)=>data_re_out(1703),
            data_re_out(54)=>data_re_out(1735),
            data_re_out(55)=>data_re_out(1767),
            data_re_out(56)=>data_re_out(1799),
            data_re_out(57)=>data_re_out(1831),
            data_re_out(58)=>data_re_out(1863),
            data_re_out(59)=>data_re_out(1895),
            data_re_out(60)=>data_re_out(1927),
            data_re_out(61)=>data_re_out(1959),
            data_re_out(62)=>data_re_out(1991),
            data_re_out(63)=>data_re_out(2023),
            data_im_out(0)=>data_im_out(7),
            data_im_out(1)=>data_im_out(39),
            data_im_out(2)=>data_im_out(71),
            data_im_out(3)=>data_im_out(103),
            data_im_out(4)=>data_im_out(135),
            data_im_out(5)=>data_im_out(167),
            data_im_out(6)=>data_im_out(199),
            data_im_out(7)=>data_im_out(231),
            data_im_out(8)=>data_im_out(263),
            data_im_out(9)=>data_im_out(295),
            data_im_out(10)=>data_im_out(327),
            data_im_out(11)=>data_im_out(359),
            data_im_out(12)=>data_im_out(391),
            data_im_out(13)=>data_im_out(423),
            data_im_out(14)=>data_im_out(455),
            data_im_out(15)=>data_im_out(487),
            data_im_out(16)=>data_im_out(519),
            data_im_out(17)=>data_im_out(551),
            data_im_out(18)=>data_im_out(583),
            data_im_out(19)=>data_im_out(615),
            data_im_out(20)=>data_im_out(647),
            data_im_out(21)=>data_im_out(679),
            data_im_out(22)=>data_im_out(711),
            data_im_out(23)=>data_im_out(743),
            data_im_out(24)=>data_im_out(775),
            data_im_out(25)=>data_im_out(807),
            data_im_out(26)=>data_im_out(839),
            data_im_out(27)=>data_im_out(871),
            data_im_out(28)=>data_im_out(903),
            data_im_out(29)=>data_im_out(935),
            data_im_out(30)=>data_im_out(967),
            data_im_out(31)=>data_im_out(999),
            data_im_out(32)=>data_im_out(1031),
            data_im_out(33)=>data_im_out(1063),
            data_im_out(34)=>data_im_out(1095),
            data_im_out(35)=>data_im_out(1127),
            data_im_out(36)=>data_im_out(1159),
            data_im_out(37)=>data_im_out(1191),
            data_im_out(38)=>data_im_out(1223),
            data_im_out(39)=>data_im_out(1255),
            data_im_out(40)=>data_im_out(1287),
            data_im_out(41)=>data_im_out(1319),
            data_im_out(42)=>data_im_out(1351),
            data_im_out(43)=>data_im_out(1383),
            data_im_out(44)=>data_im_out(1415),
            data_im_out(45)=>data_im_out(1447),
            data_im_out(46)=>data_im_out(1479),
            data_im_out(47)=>data_im_out(1511),
            data_im_out(48)=>data_im_out(1543),
            data_im_out(49)=>data_im_out(1575),
            data_im_out(50)=>data_im_out(1607),
            data_im_out(51)=>data_im_out(1639),
            data_im_out(52)=>data_im_out(1671),
            data_im_out(53)=>data_im_out(1703),
            data_im_out(54)=>data_im_out(1735),
            data_im_out(55)=>data_im_out(1767),
            data_im_out(56)=>data_im_out(1799),
            data_im_out(57)=>data_im_out(1831),
            data_im_out(58)=>data_im_out(1863),
            data_im_out(59)=>data_im_out(1895),
            data_im_out(60)=>data_im_out(1927),
            data_im_out(61)=>data_im_out(1959),
            data_im_out(62)=>data_im_out(1991),
            data_im_out(63)=>data_im_out(2023)
        );           

    URFFT_PT64_8 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(8),
            data_re_in(1)=>mul_re_out(40),
            data_re_in(2)=>mul_re_out(72),
            data_re_in(3)=>mul_re_out(104),
            data_re_in(4)=>mul_re_out(136),
            data_re_in(5)=>mul_re_out(168),
            data_re_in(6)=>mul_re_out(200),
            data_re_in(7)=>mul_re_out(232),
            data_re_in(8)=>mul_re_out(264),
            data_re_in(9)=>mul_re_out(296),
            data_re_in(10)=>mul_re_out(328),
            data_re_in(11)=>mul_re_out(360),
            data_re_in(12)=>mul_re_out(392),
            data_re_in(13)=>mul_re_out(424),
            data_re_in(14)=>mul_re_out(456),
            data_re_in(15)=>mul_re_out(488),
            data_re_in(16)=>mul_re_out(520),
            data_re_in(17)=>mul_re_out(552),
            data_re_in(18)=>mul_re_out(584),
            data_re_in(19)=>mul_re_out(616),
            data_re_in(20)=>mul_re_out(648),
            data_re_in(21)=>mul_re_out(680),
            data_re_in(22)=>mul_re_out(712),
            data_re_in(23)=>mul_re_out(744),
            data_re_in(24)=>mul_re_out(776),
            data_re_in(25)=>mul_re_out(808),
            data_re_in(26)=>mul_re_out(840),
            data_re_in(27)=>mul_re_out(872),
            data_re_in(28)=>mul_re_out(904),
            data_re_in(29)=>mul_re_out(936),
            data_re_in(30)=>mul_re_out(968),
            data_re_in(31)=>mul_re_out(1000),
            data_re_in(32)=>mul_re_out(1032),
            data_re_in(33)=>mul_re_out(1064),
            data_re_in(34)=>mul_re_out(1096),
            data_re_in(35)=>mul_re_out(1128),
            data_re_in(36)=>mul_re_out(1160),
            data_re_in(37)=>mul_re_out(1192),
            data_re_in(38)=>mul_re_out(1224),
            data_re_in(39)=>mul_re_out(1256),
            data_re_in(40)=>mul_re_out(1288),
            data_re_in(41)=>mul_re_out(1320),
            data_re_in(42)=>mul_re_out(1352),
            data_re_in(43)=>mul_re_out(1384),
            data_re_in(44)=>mul_re_out(1416),
            data_re_in(45)=>mul_re_out(1448),
            data_re_in(46)=>mul_re_out(1480),
            data_re_in(47)=>mul_re_out(1512),
            data_re_in(48)=>mul_re_out(1544),
            data_re_in(49)=>mul_re_out(1576),
            data_re_in(50)=>mul_re_out(1608),
            data_re_in(51)=>mul_re_out(1640),
            data_re_in(52)=>mul_re_out(1672),
            data_re_in(53)=>mul_re_out(1704),
            data_re_in(54)=>mul_re_out(1736),
            data_re_in(55)=>mul_re_out(1768),
            data_re_in(56)=>mul_re_out(1800),
            data_re_in(57)=>mul_re_out(1832),
            data_re_in(58)=>mul_re_out(1864),
            data_re_in(59)=>mul_re_out(1896),
            data_re_in(60)=>mul_re_out(1928),
            data_re_in(61)=>mul_re_out(1960),
            data_re_in(62)=>mul_re_out(1992),
            data_re_in(63)=>mul_re_out(2024),
            data_im_in(0)=>mul_im_out(8),
            data_im_in(1)=>mul_im_out(40),
            data_im_in(2)=>mul_im_out(72),
            data_im_in(3)=>mul_im_out(104),
            data_im_in(4)=>mul_im_out(136),
            data_im_in(5)=>mul_im_out(168),
            data_im_in(6)=>mul_im_out(200),
            data_im_in(7)=>mul_im_out(232),
            data_im_in(8)=>mul_im_out(264),
            data_im_in(9)=>mul_im_out(296),
            data_im_in(10)=>mul_im_out(328),
            data_im_in(11)=>mul_im_out(360),
            data_im_in(12)=>mul_im_out(392),
            data_im_in(13)=>mul_im_out(424),
            data_im_in(14)=>mul_im_out(456),
            data_im_in(15)=>mul_im_out(488),
            data_im_in(16)=>mul_im_out(520),
            data_im_in(17)=>mul_im_out(552),
            data_im_in(18)=>mul_im_out(584),
            data_im_in(19)=>mul_im_out(616),
            data_im_in(20)=>mul_im_out(648),
            data_im_in(21)=>mul_im_out(680),
            data_im_in(22)=>mul_im_out(712),
            data_im_in(23)=>mul_im_out(744),
            data_im_in(24)=>mul_im_out(776),
            data_im_in(25)=>mul_im_out(808),
            data_im_in(26)=>mul_im_out(840),
            data_im_in(27)=>mul_im_out(872),
            data_im_in(28)=>mul_im_out(904),
            data_im_in(29)=>mul_im_out(936),
            data_im_in(30)=>mul_im_out(968),
            data_im_in(31)=>mul_im_out(1000),
            data_im_in(32)=>mul_im_out(1032),
            data_im_in(33)=>mul_im_out(1064),
            data_im_in(34)=>mul_im_out(1096),
            data_im_in(35)=>mul_im_out(1128),
            data_im_in(36)=>mul_im_out(1160),
            data_im_in(37)=>mul_im_out(1192),
            data_im_in(38)=>mul_im_out(1224),
            data_im_in(39)=>mul_im_out(1256),
            data_im_in(40)=>mul_im_out(1288),
            data_im_in(41)=>mul_im_out(1320),
            data_im_in(42)=>mul_im_out(1352),
            data_im_in(43)=>mul_im_out(1384),
            data_im_in(44)=>mul_im_out(1416),
            data_im_in(45)=>mul_im_out(1448),
            data_im_in(46)=>mul_im_out(1480),
            data_im_in(47)=>mul_im_out(1512),
            data_im_in(48)=>mul_im_out(1544),
            data_im_in(49)=>mul_im_out(1576),
            data_im_in(50)=>mul_im_out(1608),
            data_im_in(51)=>mul_im_out(1640),
            data_im_in(52)=>mul_im_out(1672),
            data_im_in(53)=>mul_im_out(1704),
            data_im_in(54)=>mul_im_out(1736),
            data_im_in(55)=>mul_im_out(1768),
            data_im_in(56)=>mul_im_out(1800),
            data_im_in(57)=>mul_im_out(1832),
            data_im_in(58)=>mul_im_out(1864),
            data_im_in(59)=>mul_im_out(1896),
            data_im_in(60)=>mul_im_out(1928),
            data_im_in(61)=>mul_im_out(1960),
            data_im_in(62)=>mul_im_out(1992),
            data_im_in(63)=>mul_im_out(2024),
            data_re_out(0)=>data_re_out(8),
            data_re_out(1)=>data_re_out(40),
            data_re_out(2)=>data_re_out(72),
            data_re_out(3)=>data_re_out(104),
            data_re_out(4)=>data_re_out(136),
            data_re_out(5)=>data_re_out(168),
            data_re_out(6)=>data_re_out(200),
            data_re_out(7)=>data_re_out(232),
            data_re_out(8)=>data_re_out(264),
            data_re_out(9)=>data_re_out(296),
            data_re_out(10)=>data_re_out(328),
            data_re_out(11)=>data_re_out(360),
            data_re_out(12)=>data_re_out(392),
            data_re_out(13)=>data_re_out(424),
            data_re_out(14)=>data_re_out(456),
            data_re_out(15)=>data_re_out(488),
            data_re_out(16)=>data_re_out(520),
            data_re_out(17)=>data_re_out(552),
            data_re_out(18)=>data_re_out(584),
            data_re_out(19)=>data_re_out(616),
            data_re_out(20)=>data_re_out(648),
            data_re_out(21)=>data_re_out(680),
            data_re_out(22)=>data_re_out(712),
            data_re_out(23)=>data_re_out(744),
            data_re_out(24)=>data_re_out(776),
            data_re_out(25)=>data_re_out(808),
            data_re_out(26)=>data_re_out(840),
            data_re_out(27)=>data_re_out(872),
            data_re_out(28)=>data_re_out(904),
            data_re_out(29)=>data_re_out(936),
            data_re_out(30)=>data_re_out(968),
            data_re_out(31)=>data_re_out(1000),
            data_re_out(32)=>data_re_out(1032),
            data_re_out(33)=>data_re_out(1064),
            data_re_out(34)=>data_re_out(1096),
            data_re_out(35)=>data_re_out(1128),
            data_re_out(36)=>data_re_out(1160),
            data_re_out(37)=>data_re_out(1192),
            data_re_out(38)=>data_re_out(1224),
            data_re_out(39)=>data_re_out(1256),
            data_re_out(40)=>data_re_out(1288),
            data_re_out(41)=>data_re_out(1320),
            data_re_out(42)=>data_re_out(1352),
            data_re_out(43)=>data_re_out(1384),
            data_re_out(44)=>data_re_out(1416),
            data_re_out(45)=>data_re_out(1448),
            data_re_out(46)=>data_re_out(1480),
            data_re_out(47)=>data_re_out(1512),
            data_re_out(48)=>data_re_out(1544),
            data_re_out(49)=>data_re_out(1576),
            data_re_out(50)=>data_re_out(1608),
            data_re_out(51)=>data_re_out(1640),
            data_re_out(52)=>data_re_out(1672),
            data_re_out(53)=>data_re_out(1704),
            data_re_out(54)=>data_re_out(1736),
            data_re_out(55)=>data_re_out(1768),
            data_re_out(56)=>data_re_out(1800),
            data_re_out(57)=>data_re_out(1832),
            data_re_out(58)=>data_re_out(1864),
            data_re_out(59)=>data_re_out(1896),
            data_re_out(60)=>data_re_out(1928),
            data_re_out(61)=>data_re_out(1960),
            data_re_out(62)=>data_re_out(1992),
            data_re_out(63)=>data_re_out(2024),
            data_im_out(0)=>data_im_out(8),
            data_im_out(1)=>data_im_out(40),
            data_im_out(2)=>data_im_out(72),
            data_im_out(3)=>data_im_out(104),
            data_im_out(4)=>data_im_out(136),
            data_im_out(5)=>data_im_out(168),
            data_im_out(6)=>data_im_out(200),
            data_im_out(7)=>data_im_out(232),
            data_im_out(8)=>data_im_out(264),
            data_im_out(9)=>data_im_out(296),
            data_im_out(10)=>data_im_out(328),
            data_im_out(11)=>data_im_out(360),
            data_im_out(12)=>data_im_out(392),
            data_im_out(13)=>data_im_out(424),
            data_im_out(14)=>data_im_out(456),
            data_im_out(15)=>data_im_out(488),
            data_im_out(16)=>data_im_out(520),
            data_im_out(17)=>data_im_out(552),
            data_im_out(18)=>data_im_out(584),
            data_im_out(19)=>data_im_out(616),
            data_im_out(20)=>data_im_out(648),
            data_im_out(21)=>data_im_out(680),
            data_im_out(22)=>data_im_out(712),
            data_im_out(23)=>data_im_out(744),
            data_im_out(24)=>data_im_out(776),
            data_im_out(25)=>data_im_out(808),
            data_im_out(26)=>data_im_out(840),
            data_im_out(27)=>data_im_out(872),
            data_im_out(28)=>data_im_out(904),
            data_im_out(29)=>data_im_out(936),
            data_im_out(30)=>data_im_out(968),
            data_im_out(31)=>data_im_out(1000),
            data_im_out(32)=>data_im_out(1032),
            data_im_out(33)=>data_im_out(1064),
            data_im_out(34)=>data_im_out(1096),
            data_im_out(35)=>data_im_out(1128),
            data_im_out(36)=>data_im_out(1160),
            data_im_out(37)=>data_im_out(1192),
            data_im_out(38)=>data_im_out(1224),
            data_im_out(39)=>data_im_out(1256),
            data_im_out(40)=>data_im_out(1288),
            data_im_out(41)=>data_im_out(1320),
            data_im_out(42)=>data_im_out(1352),
            data_im_out(43)=>data_im_out(1384),
            data_im_out(44)=>data_im_out(1416),
            data_im_out(45)=>data_im_out(1448),
            data_im_out(46)=>data_im_out(1480),
            data_im_out(47)=>data_im_out(1512),
            data_im_out(48)=>data_im_out(1544),
            data_im_out(49)=>data_im_out(1576),
            data_im_out(50)=>data_im_out(1608),
            data_im_out(51)=>data_im_out(1640),
            data_im_out(52)=>data_im_out(1672),
            data_im_out(53)=>data_im_out(1704),
            data_im_out(54)=>data_im_out(1736),
            data_im_out(55)=>data_im_out(1768),
            data_im_out(56)=>data_im_out(1800),
            data_im_out(57)=>data_im_out(1832),
            data_im_out(58)=>data_im_out(1864),
            data_im_out(59)=>data_im_out(1896),
            data_im_out(60)=>data_im_out(1928),
            data_im_out(61)=>data_im_out(1960),
            data_im_out(62)=>data_im_out(1992),
            data_im_out(63)=>data_im_out(2024)
        );           

    URFFT_PT64_9 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(9),
            data_re_in(1)=>mul_re_out(41),
            data_re_in(2)=>mul_re_out(73),
            data_re_in(3)=>mul_re_out(105),
            data_re_in(4)=>mul_re_out(137),
            data_re_in(5)=>mul_re_out(169),
            data_re_in(6)=>mul_re_out(201),
            data_re_in(7)=>mul_re_out(233),
            data_re_in(8)=>mul_re_out(265),
            data_re_in(9)=>mul_re_out(297),
            data_re_in(10)=>mul_re_out(329),
            data_re_in(11)=>mul_re_out(361),
            data_re_in(12)=>mul_re_out(393),
            data_re_in(13)=>mul_re_out(425),
            data_re_in(14)=>mul_re_out(457),
            data_re_in(15)=>mul_re_out(489),
            data_re_in(16)=>mul_re_out(521),
            data_re_in(17)=>mul_re_out(553),
            data_re_in(18)=>mul_re_out(585),
            data_re_in(19)=>mul_re_out(617),
            data_re_in(20)=>mul_re_out(649),
            data_re_in(21)=>mul_re_out(681),
            data_re_in(22)=>mul_re_out(713),
            data_re_in(23)=>mul_re_out(745),
            data_re_in(24)=>mul_re_out(777),
            data_re_in(25)=>mul_re_out(809),
            data_re_in(26)=>mul_re_out(841),
            data_re_in(27)=>mul_re_out(873),
            data_re_in(28)=>mul_re_out(905),
            data_re_in(29)=>mul_re_out(937),
            data_re_in(30)=>mul_re_out(969),
            data_re_in(31)=>mul_re_out(1001),
            data_re_in(32)=>mul_re_out(1033),
            data_re_in(33)=>mul_re_out(1065),
            data_re_in(34)=>mul_re_out(1097),
            data_re_in(35)=>mul_re_out(1129),
            data_re_in(36)=>mul_re_out(1161),
            data_re_in(37)=>mul_re_out(1193),
            data_re_in(38)=>mul_re_out(1225),
            data_re_in(39)=>mul_re_out(1257),
            data_re_in(40)=>mul_re_out(1289),
            data_re_in(41)=>mul_re_out(1321),
            data_re_in(42)=>mul_re_out(1353),
            data_re_in(43)=>mul_re_out(1385),
            data_re_in(44)=>mul_re_out(1417),
            data_re_in(45)=>mul_re_out(1449),
            data_re_in(46)=>mul_re_out(1481),
            data_re_in(47)=>mul_re_out(1513),
            data_re_in(48)=>mul_re_out(1545),
            data_re_in(49)=>mul_re_out(1577),
            data_re_in(50)=>mul_re_out(1609),
            data_re_in(51)=>mul_re_out(1641),
            data_re_in(52)=>mul_re_out(1673),
            data_re_in(53)=>mul_re_out(1705),
            data_re_in(54)=>mul_re_out(1737),
            data_re_in(55)=>mul_re_out(1769),
            data_re_in(56)=>mul_re_out(1801),
            data_re_in(57)=>mul_re_out(1833),
            data_re_in(58)=>mul_re_out(1865),
            data_re_in(59)=>mul_re_out(1897),
            data_re_in(60)=>mul_re_out(1929),
            data_re_in(61)=>mul_re_out(1961),
            data_re_in(62)=>mul_re_out(1993),
            data_re_in(63)=>mul_re_out(2025),
            data_im_in(0)=>mul_im_out(9),
            data_im_in(1)=>mul_im_out(41),
            data_im_in(2)=>mul_im_out(73),
            data_im_in(3)=>mul_im_out(105),
            data_im_in(4)=>mul_im_out(137),
            data_im_in(5)=>mul_im_out(169),
            data_im_in(6)=>mul_im_out(201),
            data_im_in(7)=>mul_im_out(233),
            data_im_in(8)=>mul_im_out(265),
            data_im_in(9)=>mul_im_out(297),
            data_im_in(10)=>mul_im_out(329),
            data_im_in(11)=>mul_im_out(361),
            data_im_in(12)=>mul_im_out(393),
            data_im_in(13)=>mul_im_out(425),
            data_im_in(14)=>mul_im_out(457),
            data_im_in(15)=>mul_im_out(489),
            data_im_in(16)=>mul_im_out(521),
            data_im_in(17)=>mul_im_out(553),
            data_im_in(18)=>mul_im_out(585),
            data_im_in(19)=>mul_im_out(617),
            data_im_in(20)=>mul_im_out(649),
            data_im_in(21)=>mul_im_out(681),
            data_im_in(22)=>mul_im_out(713),
            data_im_in(23)=>mul_im_out(745),
            data_im_in(24)=>mul_im_out(777),
            data_im_in(25)=>mul_im_out(809),
            data_im_in(26)=>mul_im_out(841),
            data_im_in(27)=>mul_im_out(873),
            data_im_in(28)=>mul_im_out(905),
            data_im_in(29)=>mul_im_out(937),
            data_im_in(30)=>mul_im_out(969),
            data_im_in(31)=>mul_im_out(1001),
            data_im_in(32)=>mul_im_out(1033),
            data_im_in(33)=>mul_im_out(1065),
            data_im_in(34)=>mul_im_out(1097),
            data_im_in(35)=>mul_im_out(1129),
            data_im_in(36)=>mul_im_out(1161),
            data_im_in(37)=>mul_im_out(1193),
            data_im_in(38)=>mul_im_out(1225),
            data_im_in(39)=>mul_im_out(1257),
            data_im_in(40)=>mul_im_out(1289),
            data_im_in(41)=>mul_im_out(1321),
            data_im_in(42)=>mul_im_out(1353),
            data_im_in(43)=>mul_im_out(1385),
            data_im_in(44)=>mul_im_out(1417),
            data_im_in(45)=>mul_im_out(1449),
            data_im_in(46)=>mul_im_out(1481),
            data_im_in(47)=>mul_im_out(1513),
            data_im_in(48)=>mul_im_out(1545),
            data_im_in(49)=>mul_im_out(1577),
            data_im_in(50)=>mul_im_out(1609),
            data_im_in(51)=>mul_im_out(1641),
            data_im_in(52)=>mul_im_out(1673),
            data_im_in(53)=>mul_im_out(1705),
            data_im_in(54)=>mul_im_out(1737),
            data_im_in(55)=>mul_im_out(1769),
            data_im_in(56)=>mul_im_out(1801),
            data_im_in(57)=>mul_im_out(1833),
            data_im_in(58)=>mul_im_out(1865),
            data_im_in(59)=>mul_im_out(1897),
            data_im_in(60)=>mul_im_out(1929),
            data_im_in(61)=>mul_im_out(1961),
            data_im_in(62)=>mul_im_out(1993),
            data_im_in(63)=>mul_im_out(2025),
            data_re_out(0)=>data_re_out(9),
            data_re_out(1)=>data_re_out(41),
            data_re_out(2)=>data_re_out(73),
            data_re_out(3)=>data_re_out(105),
            data_re_out(4)=>data_re_out(137),
            data_re_out(5)=>data_re_out(169),
            data_re_out(6)=>data_re_out(201),
            data_re_out(7)=>data_re_out(233),
            data_re_out(8)=>data_re_out(265),
            data_re_out(9)=>data_re_out(297),
            data_re_out(10)=>data_re_out(329),
            data_re_out(11)=>data_re_out(361),
            data_re_out(12)=>data_re_out(393),
            data_re_out(13)=>data_re_out(425),
            data_re_out(14)=>data_re_out(457),
            data_re_out(15)=>data_re_out(489),
            data_re_out(16)=>data_re_out(521),
            data_re_out(17)=>data_re_out(553),
            data_re_out(18)=>data_re_out(585),
            data_re_out(19)=>data_re_out(617),
            data_re_out(20)=>data_re_out(649),
            data_re_out(21)=>data_re_out(681),
            data_re_out(22)=>data_re_out(713),
            data_re_out(23)=>data_re_out(745),
            data_re_out(24)=>data_re_out(777),
            data_re_out(25)=>data_re_out(809),
            data_re_out(26)=>data_re_out(841),
            data_re_out(27)=>data_re_out(873),
            data_re_out(28)=>data_re_out(905),
            data_re_out(29)=>data_re_out(937),
            data_re_out(30)=>data_re_out(969),
            data_re_out(31)=>data_re_out(1001),
            data_re_out(32)=>data_re_out(1033),
            data_re_out(33)=>data_re_out(1065),
            data_re_out(34)=>data_re_out(1097),
            data_re_out(35)=>data_re_out(1129),
            data_re_out(36)=>data_re_out(1161),
            data_re_out(37)=>data_re_out(1193),
            data_re_out(38)=>data_re_out(1225),
            data_re_out(39)=>data_re_out(1257),
            data_re_out(40)=>data_re_out(1289),
            data_re_out(41)=>data_re_out(1321),
            data_re_out(42)=>data_re_out(1353),
            data_re_out(43)=>data_re_out(1385),
            data_re_out(44)=>data_re_out(1417),
            data_re_out(45)=>data_re_out(1449),
            data_re_out(46)=>data_re_out(1481),
            data_re_out(47)=>data_re_out(1513),
            data_re_out(48)=>data_re_out(1545),
            data_re_out(49)=>data_re_out(1577),
            data_re_out(50)=>data_re_out(1609),
            data_re_out(51)=>data_re_out(1641),
            data_re_out(52)=>data_re_out(1673),
            data_re_out(53)=>data_re_out(1705),
            data_re_out(54)=>data_re_out(1737),
            data_re_out(55)=>data_re_out(1769),
            data_re_out(56)=>data_re_out(1801),
            data_re_out(57)=>data_re_out(1833),
            data_re_out(58)=>data_re_out(1865),
            data_re_out(59)=>data_re_out(1897),
            data_re_out(60)=>data_re_out(1929),
            data_re_out(61)=>data_re_out(1961),
            data_re_out(62)=>data_re_out(1993),
            data_re_out(63)=>data_re_out(2025),
            data_im_out(0)=>data_im_out(9),
            data_im_out(1)=>data_im_out(41),
            data_im_out(2)=>data_im_out(73),
            data_im_out(3)=>data_im_out(105),
            data_im_out(4)=>data_im_out(137),
            data_im_out(5)=>data_im_out(169),
            data_im_out(6)=>data_im_out(201),
            data_im_out(7)=>data_im_out(233),
            data_im_out(8)=>data_im_out(265),
            data_im_out(9)=>data_im_out(297),
            data_im_out(10)=>data_im_out(329),
            data_im_out(11)=>data_im_out(361),
            data_im_out(12)=>data_im_out(393),
            data_im_out(13)=>data_im_out(425),
            data_im_out(14)=>data_im_out(457),
            data_im_out(15)=>data_im_out(489),
            data_im_out(16)=>data_im_out(521),
            data_im_out(17)=>data_im_out(553),
            data_im_out(18)=>data_im_out(585),
            data_im_out(19)=>data_im_out(617),
            data_im_out(20)=>data_im_out(649),
            data_im_out(21)=>data_im_out(681),
            data_im_out(22)=>data_im_out(713),
            data_im_out(23)=>data_im_out(745),
            data_im_out(24)=>data_im_out(777),
            data_im_out(25)=>data_im_out(809),
            data_im_out(26)=>data_im_out(841),
            data_im_out(27)=>data_im_out(873),
            data_im_out(28)=>data_im_out(905),
            data_im_out(29)=>data_im_out(937),
            data_im_out(30)=>data_im_out(969),
            data_im_out(31)=>data_im_out(1001),
            data_im_out(32)=>data_im_out(1033),
            data_im_out(33)=>data_im_out(1065),
            data_im_out(34)=>data_im_out(1097),
            data_im_out(35)=>data_im_out(1129),
            data_im_out(36)=>data_im_out(1161),
            data_im_out(37)=>data_im_out(1193),
            data_im_out(38)=>data_im_out(1225),
            data_im_out(39)=>data_im_out(1257),
            data_im_out(40)=>data_im_out(1289),
            data_im_out(41)=>data_im_out(1321),
            data_im_out(42)=>data_im_out(1353),
            data_im_out(43)=>data_im_out(1385),
            data_im_out(44)=>data_im_out(1417),
            data_im_out(45)=>data_im_out(1449),
            data_im_out(46)=>data_im_out(1481),
            data_im_out(47)=>data_im_out(1513),
            data_im_out(48)=>data_im_out(1545),
            data_im_out(49)=>data_im_out(1577),
            data_im_out(50)=>data_im_out(1609),
            data_im_out(51)=>data_im_out(1641),
            data_im_out(52)=>data_im_out(1673),
            data_im_out(53)=>data_im_out(1705),
            data_im_out(54)=>data_im_out(1737),
            data_im_out(55)=>data_im_out(1769),
            data_im_out(56)=>data_im_out(1801),
            data_im_out(57)=>data_im_out(1833),
            data_im_out(58)=>data_im_out(1865),
            data_im_out(59)=>data_im_out(1897),
            data_im_out(60)=>data_im_out(1929),
            data_im_out(61)=>data_im_out(1961),
            data_im_out(62)=>data_im_out(1993),
            data_im_out(63)=>data_im_out(2025)
        );           

    URFFT_PT64_10 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(10),
            data_re_in(1)=>mul_re_out(42),
            data_re_in(2)=>mul_re_out(74),
            data_re_in(3)=>mul_re_out(106),
            data_re_in(4)=>mul_re_out(138),
            data_re_in(5)=>mul_re_out(170),
            data_re_in(6)=>mul_re_out(202),
            data_re_in(7)=>mul_re_out(234),
            data_re_in(8)=>mul_re_out(266),
            data_re_in(9)=>mul_re_out(298),
            data_re_in(10)=>mul_re_out(330),
            data_re_in(11)=>mul_re_out(362),
            data_re_in(12)=>mul_re_out(394),
            data_re_in(13)=>mul_re_out(426),
            data_re_in(14)=>mul_re_out(458),
            data_re_in(15)=>mul_re_out(490),
            data_re_in(16)=>mul_re_out(522),
            data_re_in(17)=>mul_re_out(554),
            data_re_in(18)=>mul_re_out(586),
            data_re_in(19)=>mul_re_out(618),
            data_re_in(20)=>mul_re_out(650),
            data_re_in(21)=>mul_re_out(682),
            data_re_in(22)=>mul_re_out(714),
            data_re_in(23)=>mul_re_out(746),
            data_re_in(24)=>mul_re_out(778),
            data_re_in(25)=>mul_re_out(810),
            data_re_in(26)=>mul_re_out(842),
            data_re_in(27)=>mul_re_out(874),
            data_re_in(28)=>mul_re_out(906),
            data_re_in(29)=>mul_re_out(938),
            data_re_in(30)=>mul_re_out(970),
            data_re_in(31)=>mul_re_out(1002),
            data_re_in(32)=>mul_re_out(1034),
            data_re_in(33)=>mul_re_out(1066),
            data_re_in(34)=>mul_re_out(1098),
            data_re_in(35)=>mul_re_out(1130),
            data_re_in(36)=>mul_re_out(1162),
            data_re_in(37)=>mul_re_out(1194),
            data_re_in(38)=>mul_re_out(1226),
            data_re_in(39)=>mul_re_out(1258),
            data_re_in(40)=>mul_re_out(1290),
            data_re_in(41)=>mul_re_out(1322),
            data_re_in(42)=>mul_re_out(1354),
            data_re_in(43)=>mul_re_out(1386),
            data_re_in(44)=>mul_re_out(1418),
            data_re_in(45)=>mul_re_out(1450),
            data_re_in(46)=>mul_re_out(1482),
            data_re_in(47)=>mul_re_out(1514),
            data_re_in(48)=>mul_re_out(1546),
            data_re_in(49)=>mul_re_out(1578),
            data_re_in(50)=>mul_re_out(1610),
            data_re_in(51)=>mul_re_out(1642),
            data_re_in(52)=>mul_re_out(1674),
            data_re_in(53)=>mul_re_out(1706),
            data_re_in(54)=>mul_re_out(1738),
            data_re_in(55)=>mul_re_out(1770),
            data_re_in(56)=>mul_re_out(1802),
            data_re_in(57)=>mul_re_out(1834),
            data_re_in(58)=>mul_re_out(1866),
            data_re_in(59)=>mul_re_out(1898),
            data_re_in(60)=>mul_re_out(1930),
            data_re_in(61)=>mul_re_out(1962),
            data_re_in(62)=>mul_re_out(1994),
            data_re_in(63)=>mul_re_out(2026),
            data_im_in(0)=>mul_im_out(10),
            data_im_in(1)=>mul_im_out(42),
            data_im_in(2)=>mul_im_out(74),
            data_im_in(3)=>mul_im_out(106),
            data_im_in(4)=>mul_im_out(138),
            data_im_in(5)=>mul_im_out(170),
            data_im_in(6)=>mul_im_out(202),
            data_im_in(7)=>mul_im_out(234),
            data_im_in(8)=>mul_im_out(266),
            data_im_in(9)=>mul_im_out(298),
            data_im_in(10)=>mul_im_out(330),
            data_im_in(11)=>mul_im_out(362),
            data_im_in(12)=>mul_im_out(394),
            data_im_in(13)=>mul_im_out(426),
            data_im_in(14)=>mul_im_out(458),
            data_im_in(15)=>mul_im_out(490),
            data_im_in(16)=>mul_im_out(522),
            data_im_in(17)=>mul_im_out(554),
            data_im_in(18)=>mul_im_out(586),
            data_im_in(19)=>mul_im_out(618),
            data_im_in(20)=>mul_im_out(650),
            data_im_in(21)=>mul_im_out(682),
            data_im_in(22)=>mul_im_out(714),
            data_im_in(23)=>mul_im_out(746),
            data_im_in(24)=>mul_im_out(778),
            data_im_in(25)=>mul_im_out(810),
            data_im_in(26)=>mul_im_out(842),
            data_im_in(27)=>mul_im_out(874),
            data_im_in(28)=>mul_im_out(906),
            data_im_in(29)=>mul_im_out(938),
            data_im_in(30)=>mul_im_out(970),
            data_im_in(31)=>mul_im_out(1002),
            data_im_in(32)=>mul_im_out(1034),
            data_im_in(33)=>mul_im_out(1066),
            data_im_in(34)=>mul_im_out(1098),
            data_im_in(35)=>mul_im_out(1130),
            data_im_in(36)=>mul_im_out(1162),
            data_im_in(37)=>mul_im_out(1194),
            data_im_in(38)=>mul_im_out(1226),
            data_im_in(39)=>mul_im_out(1258),
            data_im_in(40)=>mul_im_out(1290),
            data_im_in(41)=>mul_im_out(1322),
            data_im_in(42)=>mul_im_out(1354),
            data_im_in(43)=>mul_im_out(1386),
            data_im_in(44)=>mul_im_out(1418),
            data_im_in(45)=>mul_im_out(1450),
            data_im_in(46)=>mul_im_out(1482),
            data_im_in(47)=>mul_im_out(1514),
            data_im_in(48)=>mul_im_out(1546),
            data_im_in(49)=>mul_im_out(1578),
            data_im_in(50)=>mul_im_out(1610),
            data_im_in(51)=>mul_im_out(1642),
            data_im_in(52)=>mul_im_out(1674),
            data_im_in(53)=>mul_im_out(1706),
            data_im_in(54)=>mul_im_out(1738),
            data_im_in(55)=>mul_im_out(1770),
            data_im_in(56)=>mul_im_out(1802),
            data_im_in(57)=>mul_im_out(1834),
            data_im_in(58)=>mul_im_out(1866),
            data_im_in(59)=>mul_im_out(1898),
            data_im_in(60)=>mul_im_out(1930),
            data_im_in(61)=>mul_im_out(1962),
            data_im_in(62)=>mul_im_out(1994),
            data_im_in(63)=>mul_im_out(2026),
            data_re_out(0)=>data_re_out(10),
            data_re_out(1)=>data_re_out(42),
            data_re_out(2)=>data_re_out(74),
            data_re_out(3)=>data_re_out(106),
            data_re_out(4)=>data_re_out(138),
            data_re_out(5)=>data_re_out(170),
            data_re_out(6)=>data_re_out(202),
            data_re_out(7)=>data_re_out(234),
            data_re_out(8)=>data_re_out(266),
            data_re_out(9)=>data_re_out(298),
            data_re_out(10)=>data_re_out(330),
            data_re_out(11)=>data_re_out(362),
            data_re_out(12)=>data_re_out(394),
            data_re_out(13)=>data_re_out(426),
            data_re_out(14)=>data_re_out(458),
            data_re_out(15)=>data_re_out(490),
            data_re_out(16)=>data_re_out(522),
            data_re_out(17)=>data_re_out(554),
            data_re_out(18)=>data_re_out(586),
            data_re_out(19)=>data_re_out(618),
            data_re_out(20)=>data_re_out(650),
            data_re_out(21)=>data_re_out(682),
            data_re_out(22)=>data_re_out(714),
            data_re_out(23)=>data_re_out(746),
            data_re_out(24)=>data_re_out(778),
            data_re_out(25)=>data_re_out(810),
            data_re_out(26)=>data_re_out(842),
            data_re_out(27)=>data_re_out(874),
            data_re_out(28)=>data_re_out(906),
            data_re_out(29)=>data_re_out(938),
            data_re_out(30)=>data_re_out(970),
            data_re_out(31)=>data_re_out(1002),
            data_re_out(32)=>data_re_out(1034),
            data_re_out(33)=>data_re_out(1066),
            data_re_out(34)=>data_re_out(1098),
            data_re_out(35)=>data_re_out(1130),
            data_re_out(36)=>data_re_out(1162),
            data_re_out(37)=>data_re_out(1194),
            data_re_out(38)=>data_re_out(1226),
            data_re_out(39)=>data_re_out(1258),
            data_re_out(40)=>data_re_out(1290),
            data_re_out(41)=>data_re_out(1322),
            data_re_out(42)=>data_re_out(1354),
            data_re_out(43)=>data_re_out(1386),
            data_re_out(44)=>data_re_out(1418),
            data_re_out(45)=>data_re_out(1450),
            data_re_out(46)=>data_re_out(1482),
            data_re_out(47)=>data_re_out(1514),
            data_re_out(48)=>data_re_out(1546),
            data_re_out(49)=>data_re_out(1578),
            data_re_out(50)=>data_re_out(1610),
            data_re_out(51)=>data_re_out(1642),
            data_re_out(52)=>data_re_out(1674),
            data_re_out(53)=>data_re_out(1706),
            data_re_out(54)=>data_re_out(1738),
            data_re_out(55)=>data_re_out(1770),
            data_re_out(56)=>data_re_out(1802),
            data_re_out(57)=>data_re_out(1834),
            data_re_out(58)=>data_re_out(1866),
            data_re_out(59)=>data_re_out(1898),
            data_re_out(60)=>data_re_out(1930),
            data_re_out(61)=>data_re_out(1962),
            data_re_out(62)=>data_re_out(1994),
            data_re_out(63)=>data_re_out(2026),
            data_im_out(0)=>data_im_out(10),
            data_im_out(1)=>data_im_out(42),
            data_im_out(2)=>data_im_out(74),
            data_im_out(3)=>data_im_out(106),
            data_im_out(4)=>data_im_out(138),
            data_im_out(5)=>data_im_out(170),
            data_im_out(6)=>data_im_out(202),
            data_im_out(7)=>data_im_out(234),
            data_im_out(8)=>data_im_out(266),
            data_im_out(9)=>data_im_out(298),
            data_im_out(10)=>data_im_out(330),
            data_im_out(11)=>data_im_out(362),
            data_im_out(12)=>data_im_out(394),
            data_im_out(13)=>data_im_out(426),
            data_im_out(14)=>data_im_out(458),
            data_im_out(15)=>data_im_out(490),
            data_im_out(16)=>data_im_out(522),
            data_im_out(17)=>data_im_out(554),
            data_im_out(18)=>data_im_out(586),
            data_im_out(19)=>data_im_out(618),
            data_im_out(20)=>data_im_out(650),
            data_im_out(21)=>data_im_out(682),
            data_im_out(22)=>data_im_out(714),
            data_im_out(23)=>data_im_out(746),
            data_im_out(24)=>data_im_out(778),
            data_im_out(25)=>data_im_out(810),
            data_im_out(26)=>data_im_out(842),
            data_im_out(27)=>data_im_out(874),
            data_im_out(28)=>data_im_out(906),
            data_im_out(29)=>data_im_out(938),
            data_im_out(30)=>data_im_out(970),
            data_im_out(31)=>data_im_out(1002),
            data_im_out(32)=>data_im_out(1034),
            data_im_out(33)=>data_im_out(1066),
            data_im_out(34)=>data_im_out(1098),
            data_im_out(35)=>data_im_out(1130),
            data_im_out(36)=>data_im_out(1162),
            data_im_out(37)=>data_im_out(1194),
            data_im_out(38)=>data_im_out(1226),
            data_im_out(39)=>data_im_out(1258),
            data_im_out(40)=>data_im_out(1290),
            data_im_out(41)=>data_im_out(1322),
            data_im_out(42)=>data_im_out(1354),
            data_im_out(43)=>data_im_out(1386),
            data_im_out(44)=>data_im_out(1418),
            data_im_out(45)=>data_im_out(1450),
            data_im_out(46)=>data_im_out(1482),
            data_im_out(47)=>data_im_out(1514),
            data_im_out(48)=>data_im_out(1546),
            data_im_out(49)=>data_im_out(1578),
            data_im_out(50)=>data_im_out(1610),
            data_im_out(51)=>data_im_out(1642),
            data_im_out(52)=>data_im_out(1674),
            data_im_out(53)=>data_im_out(1706),
            data_im_out(54)=>data_im_out(1738),
            data_im_out(55)=>data_im_out(1770),
            data_im_out(56)=>data_im_out(1802),
            data_im_out(57)=>data_im_out(1834),
            data_im_out(58)=>data_im_out(1866),
            data_im_out(59)=>data_im_out(1898),
            data_im_out(60)=>data_im_out(1930),
            data_im_out(61)=>data_im_out(1962),
            data_im_out(62)=>data_im_out(1994),
            data_im_out(63)=>data_im_out(2026)
        );           

    URFFT_PT64_11 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(11),
            data_re_in(1)=>mul_re_out(43),
            data_re_in(2)=>mul_re_out(75),
            data_re_in(3)=>mul_re_out(107),
            data_re_in(4)=>mul_re_out(139),
            data_re_in(5)=>mul_re_out(171),
            data_re_in(6)=>mul_re_out(203),
            data_re_in(7)=>mul_re_out(235),
            data_re_in(8)=>mul_re_out(267),
            data_re_in(9)=>mul_re_out(299),
            data_re_in(10)=>mul_re_out(331),
            data_re_in(11)=>mul_re_out(363),
            data_re_in(12)=>mul_re_out(395),
            data_re_in(13)=>mul_re_out(427),
            data_re_in(14)=>mul_re_out(459),
            data_re_in(15)=>mul_re_out(491),
            data_re_in(16)=>mul_re_out(523),
            data_re_in(17)=>mul_re_out(555),
            data_re_in(18)=>mul_re_out(587),
            data_re_in(19)=>mul_re_out(619),
            data_re_in(20)=>mul_re_out(651),
            data_re_in(21)=>mul_re_out(683),
            data_re_in(22)=>mul_re_out(715),
            data_re_in(23)=>mul_re_out(747),
            data_re_in(24)=>mul_re_out(779),
            data_re_in(25)=>mul_re_out(811),
            data_re_in(26)=>mul_re_out(843),
            data_re_in(27)=>mul_re_out(875),
            data_re_in(28)=>mul_re_out(907),
            data_re_in(29)=>mul_re_out(939),
            data_re_in(30)=>mul_re_out(971),
            data_re_in(31)=>mul_re_out(1003),
            data_re_in(32)=>mul_re_out(1035),
            data_re_in(33)=>mul_re_out(1067),
            data_re_in(34)=>mul_re_out(1099),
            data_re_in(35)=>mul_re_out(1131),
            data_re_in(36)=>mul_re_out(1163),
            data_re_in(37)=>mul_re_out(1195),
            data_re_in(38)=>mul_re_out(1227),
            data_re_in(39)=>mul_re_out(1259),
            data_re_in(40)=>mul_re_out(1291),
            data_re_in(41)=>mul_re_out(1323),
            data_re_in(42)=>mul_re_out(1355),
            data_re_in(43)=>mul_re_out(1387),
            data_re_in(44)=>mul_re_out(1419),
            data_re_in(45)=>mul_re_out(1451),
            data_re_in(46)=>mul_re_out(1483),
            data_re_in(47)=>mul_re_out(1515),
            data_re_in(48)=>mul_re_out(1547),
            data_re_in(49)=>mul_re_out(1579),
            data_re_in(50)=>mul_re_out(1611),
            data_re_in(51)=>mul_re_out(1643),
            data_re_in(52)=>mul_re_out(1675),
            data_re_in(53)=>mul_re_out(1707),
            data_re_in(54)=>mul_re_out(1739),
            data_re_in(55)=>mul_re_out(1771),
            data_re_in(56)=>mul_re_out(1803),
            data_re_in(57)=>mul_re_out(1835),
            data_re_in(58)=>mul_re_out(1867),
            data_re_in(59)=>mul_re_out(1899),
            data_re_in(60)=>mul_re_out(1931),
            data_re_in(61)=>mul_re_out(1963),
            data_re_in(62)=>mul_re_out(1995),
            data_re_in(63)=>mul_re_out(2027),
            data_im_in(0)=>mul_im_out(11),
            data_im_in(1)=>mul_im_out(43),
            data_im_in(2)=>mul_im_out(75),
            data_im_in(3)=>mul_im_out(107),
            data_im_in(4)=>mul_im_out(139),
            data_im_in(5)=>mul_im_out(171),
            data_im_in(6)=>mul_im_out(203),
            data_im_in(7)=>mul_im_out(235),
            data_im_in(8)=>mul_im_out(267),
            data_im_in(9)=>mul_im_out(299),
            data_im_in(10)=>mul_im_out(331),
            data_im_in(11)=>mul_im_out(363),
            data_im_in(12)=>mul_im_out(395),
            data_im_in(13)=>mul_im_out(427),
            data_im_in(14)=>mul_im_out(459),
            data_im_in(15)=>mul_im_out(491),
            data_im_in(16)=>mul_im_out(523),
            data_im_in(17)=>mul_im_out(555),
            data_im_in(18)=>mul_im_out(587),
            data_im_in(19)=>mul_im_out(619),
            data_im_in(20)=>mul_im_out(651),
            data_im_in(21)=>mul_im_out(683),
            data_im_in(22)=>mul_im_out(715),
            data_im_in(23)=>mul_im_out(747),
            data_im_in(24)=>mul_im_out(779),
            data_im_in(25)=>mul_im_out(811),
            data_im_in(26)=>mul_im_out(843),
            data_im_in(27)=>mul_im_out(875),
            data_im_in(28)=>mul_im_out(907),
            data_im_in(29)=>mul_im_out(939),
            data_im_in(30)=>mul_im_out(971),
            data_im_in(31)=>mul_im_out(1003),
            data_im_in(32)=>mul_im_out(1035),
            data_im_in(33)=>mul_im_out(1067),
            data_im_in(34)=>mul_im_out(1099),
            data_im_in(35)=>mul_im_out(1131),
            data_im_in(36)=>mul_im_out(1163),
            data_im_in(37)=>mul_im_out(1195),
            data_im_in(38)=>mul_im_out(1227),
            data_im_in(39)=>mul_im_out(1259),
            data_im_in(40)=>mul_im_out(1291),
            data_im_in(41)=>mul_im_out(1323),
            data_im_in(42)=>mul_im_out(1355),
            data_im_in(43)=>mul_im_out(1387),
            data_im_in(44)=>mul_im_out(1419),
            data_im_in(45)=>mul_im_out(1451),
            data_im_in(46)=>mul_im_out(1483),
            data_im_in(47)=>mul_im_out(1515),
            data_im_in(48)=>mul_im_out(1547),
            data_im_in(49)=>mul_im_out(1579),
            data_im_in(50)=>mul_im_out(1611),
            data_im_in(51)=>mul_im_out(1643),
            data_im_in(52)=>mul_im_out(1675),
            data_im_in(53)=>mul_im_out(1707),
            data_im_in(54)=>mul_im_out(1739),
            data_im_in(55)=>mul_im_out(1771),
            data_im_in(56)=>mul_im_out(1803),
            data_im_in(57)=>mul_im_out(1835),
            data_im_in(58)=>mul_im_out(1867),
            data_im_in(59)=>mul_im_out(1899),
            data_im_in(60)=>mul_im_out(1931),
            data_im_in(61)=>mul_im_out(1963),
            data_im_in(62)=>mul_im_out(1995),
            data_im_in(63)=>mul_im_out(2027),
            data_re_out(0)=>data_re_out(11),
            data_re_out(1)=>data_re_out(43),
            data_re_out(2)=>data_re_out(75),
            data_re_out(3)=>data_re_out(107),
            data_re_out(4)=>data_re_out(139),
            data_re_out(5)=>data_re_out(171),
            data_re_out(6)=>data_re_out(203),
            data_re_out(7)=>data_re_out(235),
            data_re_out(8)=>data_re_out(267),
            data_re_out(9)=>data_re_out(299),
            data_re_out(10)=>data_re_out(331),
            data_re_out(11)=>data_re_out(363),
            data_re_out(12)=>data_re_out(395),
            data_re_out(13)=>data_re_out(427),
            data_re_out(14)=>data_re_out(459),
            data_re_out(15)=>data_re_out(491),
            data_re_out(16)=>data_re_out(523),
            data_re_out(17)=>data_re_out(555),
            data_re_out(18)=>data_re_out(587),
            data_re_out(19)=>data_re_out(619),
            data_re_out(20)=>data_re_out(651),
            data_re_out(21)=>data_re_out(683),
            data_re_out(22)=>data_re_out(715),
            data_re_out(23)=>data_re_out(747),
            data_re_out(24)=>data_re_out(779),
            data_re_out(25)=>data_re_out(811),
            data_re_out(26)=>data_re_out(843),
            data_re_out(27)=>data_re_out(875),
            data_re_out(28)=>data_re_out(907),
            data_re_out(29)=>data_re_out(939),
            data_re_out(30)=>data_re_out(971),
            data_re_out(31)=>data_re_out(1003),
            data_re_out(32)=>data_re_out(1035),
            data_re_out(33)=>data_re_out(1067),
            data_re_out(34)=>data_re_out(1099),
            data_re_out(35)=>data_re_out(1131),
            data_re_out(36)=>data_re_out(1163),
            data_re_out(37)=>data_re_out(1195),
            data_re_out(38)=>data_re_out(1227),
            data_re_out(39)=>data_re_out(1259),
            data_re_out(40)=>data_re_out(1291),
            data_re_out(41)=>data_re_out(1323),
            data_re_out(42)=>data_re_out(1355),
            data_re_out(43)=>data_re_out(1387),
            data_re_out(44)=>data_re_out(1419),
            data_re_out(45)=>data_re_out(1451),
            data_re_out(46)=>data_re_out(1483),
            data_re_out(47)=>data_re_out(1515),
            data_re_out(48)=>data_re_out(1547),
            data_re_out(49)=>data_re_out(1579),
            data_re_out(50)=>data_re_out(1611),
            data_re_out(51)=>data_re_out(1643),
            data_re_out(52)=>data_re_out(1675),
            data_re_out(53)=>data_re_out(1707),
            data_re_out(54)=>data_re_out(1739),
            data_re_out(55)=>data_re_out(1771),
            data_re_out(56)=>data_re_out(1803),
            data_re_out(57)=>data_re_out(1835),
            data_re_out(58)=>data_re_out(1867),
            data_re_out(59)=>data_re_out(1899),
            data_re_out(60)=>data_re_out(1931),
            data_re_out(61)=>data_re_out(1963),
            data_re_out(62)=>data_re_out(1995),
            data_re_out(63)=>data_re_out(2027),
            data_im_out(0)=>data_im_out(11),
            data_im_out(1)=>data_im_out(43),
            data_im_out(2)=>data_im_out(75),
            data_im_out(3)=>data_im_out(107),
            data_im_out(4)=>data_im_out(139),
            data_im_out(5)=>data_im_out(171),
            data_im_out(6)=>data_im_out(203),
            data_im_out(7)=>data_im_out(235),
            data_im_out(8)=>data_im_out(267),
            data_im_out(9)=>data_im_out(299),
            data_im_out(10)=>data_im_out(331),
            data_im_out(11)=>data_im_out(363),
            data_im_out(12)=>data_im_out(395),
            data_im_out(13)=>data_im_out(427),
            data_im_out(14)=>data_im_out(459),
            data_im_out(15)=>data_im_out(491),
            data_im_out(16)=>data_im_out(523),
            data_im_out(17)=>data_im_out(555),
            data_im_out(18)=>data_im_out(587),
            data_im_out(19)=>data_im_out(619),
            data_im_out(20)=>data_im_out(651),
            data_im_out(21)=>data_im_out(683),
            data_im_out(22)=>data_im_out(715),
            data_im_out(23)=>data_im_out(747),
            data_im_out(24)=>data_im_out(779),
            data_im_out(25)=>data_im_out(811),
            data_im_out(26)=>data_im_out(843),
            data_im_out(27)=>data_im_out(875),
            data_im_out(28)=>data_im_out(907),
            data_im_out(29)=>data_im_out(939),
            data_im_out(30)=>data_im_out(971),
            data_im_out(31)=>data_im_out(1003),
            data_im_out(32)=>data_im_out(1035),
            data_im_out(33)=>data_im_out(1067),
            data_im_out(34)=>data_im_out(1099),
            data_im_out(35)=>data_im_out(1131),
            data_im_out(36)=>data_im_out(1163),
            data_im_out(37)=>data_im_out(1195),
            data_im_out(38)=>data_im_out(1227),
            data_im_out(39)=>data_im_out(1259),
            data_im_out(40)=>data_im_out(1291),
            data_im_out(41)=>data_im_out(1323),
            data_im_out(42)=>data_im_out(1355),
            data_im_out(43)=>data_im_out(1387),
            data_im_out(44)=>data_im_out(1419),
            data_im_out(45)=>data_im_out(1451),
            data_im_out(46)=>data_im_out(1483),
            data_im_out(47)=>data_im_out(1515),
            data_im_out(48)=>data_im_out(1547),
            data_im_out(49)=>data_im_out(1579),
            data_im_out(50)=>data_im_out(1611),
            data_im_out(51)=>data_im_out(1643),
            data_im_out(52)=>data_im_out(1675),
            data_im_out(53)=>data_im_out(1707),
            data_im_out(54)=>data_im_out(1739),
            data_im_out(55)=>data_im_out(1771),
            data_im_out(56)=>data_im_out(1803),
            data_im_out(57)=>data_im_out(1835),
            data_im_out(58)=>data_im_out(1867),
            data_im_out(59)=>data_im_out(1899),
            data_im_out(60)=>data_im_out(1931),
            data_im_out(61)=>data_im_out(1963),
            data_im_out(62)=>data_im_out(1995),
            data_im_out(63)=>data_im_out(2027)
        );           

    URFFT_PT64_12 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(12),
            data_re_in(1)=>mul_re_out(44),
            data_re_in(2)=>mul_re_out(76),
            data_re_in(3)=>mul_re_out(108),
            data_re_in(4)=>mul_re_out(140),
            data_re_in(5)=>mul_re_out(172),
            data_re_in(6)=>mul_re_out(204),
            data_re_in(7)=>mul_re_out(236),
            data_re_in(8)=>mul_re_out(268),
            data_re_in(9)=>mul_re_out(300),
            data_re_in(10)=>mul_re_out(332),
            data_re_in(11)=>mul_re_out(364),
            data_re_in(12)=>mul_re_out(396),
            data_re_in(13)=>mul_re_out(428),
            data_re_in(14)=>mul_re_out(460),
            data_re_in(15)=>mul_re_out(492),
            data_re_in(16)=>mul_re_out(524),
            data_re_in(17)=>mul_re_out(556),
            data_re_in(18)=>mul_re_out(588),
            data_re_in(19)=>mul_re_out(620),
            data_re_in(20)=>mul_re_out(652),
            data_re_in(21)=>mul_re_out(684),
            data_re_in(22)=>mul_re_out(716),
            data_re_in(23)=>mul_re_out(748),
            data_re_in(24)=>mul_re_out(780),
            data_re_in(25)=>mul_re_out(812),
            data_re_in(26)=>mul_re_out(844),
            data_re_in(27)=>mul_re_out(876),
            data_re_in(28)=>mul_re_out(908),
            data_re_in(29)=>mul_re_out(940),
            data_re_in(30)=>mul_re_out(972),
            data_re_in(31)=>mul_re_out(1004),
            data_re_in(32)=>mul_re_out(1036),
            data_re_in(33)=>mul_re_out(1068),
            data_re_in(34)=>mul_re_out(1100),
            data_re_in(35)=>mul_re_out(1132),
            data_re_in(36)=>mul_re_out(1164),
            data_re_in(37)=>mul_re_out(1196),
            data_re_in(38)=>mul_re_out(1228),
            data_re_in(39)=>mul_re_out(1260),
            data_re_in(40)=>mul_re_out(1292),
            data_re_in(41)=>mul_re_out(1324),
            data_re_in(42)=>mul_re_out(1356),
            data_re_in(43)=>mul_re_out(1388),
            data_re_in(44)=>mul_re_out(1420),
            data_re_in(45)=>mul_re_out(1452),
            data_re_in(46)=>mul_re_out(1484),
            data_re_in(47)=>mul_re_out(1516),
            data_re_in(48)=>mul_re_out(1548),
            data_re_in(49)=>mul_re_out(1580),
            data_re_in(50)=>mul_re_out(1612),
            data_re_in(51)=>mul_re_out(1644),
            data_re_in(52)=>mul_re_out(1676),
            data_re_in(53)=>mul_re_out(1708),
            data_re_in(54)=>mul_re_out(1740),
            data_re_in(55)=>mul_re_out(1772),
            data_re_in(56)=>mul_re_out(1804),
            data_re_in(57)=>mul_re_out(1836),
            data_re_in(58)=>mul_re_out(1868),
            data_re_in(59)=>mul_re_out(1900),
            data_re_in(60)=>mul_re_out(1932),
            data_re_in(61)=>mul_re_out(1964),
            data_re_in(62)=>mul_re_out(1996),
            data_re_in(63)=>mul_re_out(2028),
            data_im_in(0)=>mul_im_out(12),
            data_im_in(1)=>mul_im_out(44),
            data_im_in(2)=>mul_im_out(76),
            data_im_in(3)=>mul_im_out(108),
            data_im_in(4)=>mul_im_out(140),
            data_im_in(5)=>mul_im_out(172),
            data_im_in(6)=>mul_im_out(204),
            data_im_in(7)=>mul_im_out(236),
            data_im_in(8)=>mul_im_out(268),
            data_im_in(9)=>mul_im_out(300),
            data_im_in(10)=>mul_im_out(332),
            data_im_in(11)=>mul_im_out(364),
            data_im_in(12)=>mul_im_out(396),
            data_im_in(13)=>mul_im_out(428),
            data_im_in(14)=>mul_im_out(460),
            data_im_in(15)=>mul_im_out(492),
            data_im_in(16)=>mul_im_out(524),
            data_im_in(17)=>mul_im_out(556),
            data_im_in(18)=>mul_im_out(588),
            data_im_in(19)=>mul_im_out(620),
            data_im_in(20)=>mul_im_out(652),
            data_im_in(21)=>mul_im_out(684),
            data_im_in(22)=>mul_im_out(716),
            data_im_in(23)=>mul_im_out(748),
            data_im_in(24)=>mul_im_out(780),
            data_im_in(25)=>mul_im_out(812),
            data_im_in(26)=>mul_im_out(844),
            data_im_in(27)=>mul_im_out(876),
            data_im_in(28)=>mul_im_out(908),
            data_im_in(29)=>mul_im_out(940),
            data_im_in(30)=>mul_im_out(972),
            data_im_in(31)=>mul_im_out(1004),
            data_im_in(32)=>mul_im_out(1036),
            data_im_in(33)=>mul_im_out(1068),
            data_im_in(34)=>mul_im_out(1100),
            data_im_in(35)=>mul_im_out(1132),
            data_im_in(36)=>mul_im_out(1164),
            data_im_in(37)=>mul_im_out(1196),
            data_im_in(38)=>mul_im_out(1228),
            data_im_in(39)=>mul_im_out(1260),
            data_im_in(40)=>mul_im_out(1292),
            data_im_in(41)=>mul_im_out(1324),
            data_im_in(42)=>mul_im_out(1356),
            data_im_in(43)=>mul_im_out(1388),
            data_im_in(44)=>mul_im_out(1420),
            data_im_in(45)=>mul_im_out(1452),
            data_im_in(46)=>mul_im_out(1484),
            data_im_in(47)=>mul_im_out(1516),
            data_im_in(48)=>mul_im_out(1548),
            data_im_in(49)=>mul_im_out(1580),
            data_im_in(50)=>mul_im_out(1612),
            data_im_in(51)=>mul_im_out(1644),
            data_im_in(52)=>mul_im_out(1676),
            data_im_in(53)=>mul_im_out(1708),
            data_im_in(54)=>mul_im_out(1740),
            data_im_in(55)=>mul_im_out(1772),
            data_im_in(56)=>mul_im_out(1804),
            data_im_in(57)=>mul_im_out(1836),
            data_im_in(58)=>mul_im_out(1868),
            data_im_in(59)=>mul_im_out(1900),
            data_im_in(60)=>mul_im_out(1932),
            data_im_in(61)=>mul_im_out(1964),
            data_im_in(62)=>mul_im_out(1996),
            data_im_in(63)=>mul_im_out(2028),
            data_re_out(0)=>data_re_out(12),
            data_re_out(1)=>data_re_out(44),
            data_re_out(2)=>data_re_out(76),
            data_re_out(3)=>data_re_out(108),
            data_re_out(4)=>data_re_out(140),
            data_re_out(5)=>data_re_out(172),
            data_re_out(6)=>data_re_out(204),
            data_re_out(7)=>data_re_out(236),
            data_re_out(8)=>data_re_out(268),
            data_re_out(9)=>data_re_out(300),
            data_re_out(10)=>data_re_out(332),
            data_re_out(11)=>data_re_out(364),
            data_re_out(12)=>data_re_out(396),
            data_re_out(13)=>data_re_out(428),
            data_re_out(14)=>data_re_out(460),
            data_re_out(15)=>data_re_out(492),
            data_re_out(16)=>data_re_out(524),
            data_re_out(17)=>data_re_out(556),
            data_re_out(18)=>data_re_out(588),
            data_re_out(19)=>data_re_out(620),
            data_re_out(20)=>data_re_out(652),
            data_re_out(21)=>data_re_out(684),
            data_re_out(22)=>data_re_out(716),
            data_re_out(23)=>data_re_out(748),
            data_re_out(24)=>data_re_out(780),
            data_re_out(25)=>data_re_out(812),
            data_re_out(26)=>data_re_out(844),
            data_re_out(27)=>data_re_out(876),
            data_re_out(28)=>data_re_out(908),
            data_re_out(29)=>data_re_out(940),
            data_re_out(30)=>data_re_out(972),
            data_re_out(31)=>data_re_out(1004),
            data_re_out(32)=>data_re_out(1036),
            data_re_out(33)=>data_re_out(1068),
            data_re_out(34)=>data_re_out(1100),
            data_re_out(35)=>data_re_out(1132),
            data_re_out(36)=>data_re_out(1164),
            data_re_out(37)=>data_re_out(1196),
            data_re_out(38)=>data_re_out(1228),
            data_re_out(39)=>data_re_out(1260),
            data_re_out(40)=>data_re_out(1292),
            data_re_out(41)=>data_re_out(1324),
            data_re_out(42)=>data_re_out(1356),
            data_re_out(43)=>data_re_out(1388),
            data_re_out(44)=>data_re_out(1420),
            data_re_out(45)=>data_re_out(1452),
            data_re_out(46)=>data_re_out(1484),
            data_re_out(47)=>data_re_out(1516),
            data_re_out(48)=>data_re_out(1548),
            data_re_out(49)=>data_re_out(1580),
            data_re_out(50)=>data_re_out(1612),
            data_re_out(51)=>data_re_out(1644),
            data_re_out(52)=>data_re_out(1676),
            data_re_out(53)=>data_re_out(1708),
            data_re_out(54)=>data_re_out(1740),
            data_re_out(55)=>data_re_out(1772),
            data_re_out(56)=>data_re_out(1804),
            data_re_out(57)=>data_re_out(1836),
            data_re_out(58)=>data_re_out(1868),
            data_re_out(59)=>data_re_out(1900),
            data_re_out(60)=>data_re_out(1932),
            data_re_out(61)=>data_re_out(1964),
            data_re_out(62)=>data_re_out(1996),
            data_re_out(63)=>data_re_out(2028),
            data_im_out(0)=>data_im_out(12),
            data_im_out(1)=>data_im_out(44),
            data_im_out(2)=>data_im_out(76),
            data_im_out(3)=>data_im_out(108),
            data_im_out(4)=>data_im_out(140),
            data_im_out(5)=>data_im_out(172),
            data_im_out(6)=>data_im_out(204),
            data_im_out(7)=>data_im_out(236),
            data_im_out(8)=>data_im_out(268),
            data_im_out(9)=>data_im_out(300),
            data_im_out(10)=>data_im_out(332),
            data_im_out(11)=>data_im_out(364),
            data_im_out(12)=>data_im_out(396),
            data_im_out(13)=>data_im_out(428),
            data_im_out(14)=>data_im_out(460),
            data_im_out(15)=>data_im_out(492),
            data_im_out(16)=>data_im_out(524),
            data_im_out(17)=>data_im_out(556),
            data_im_out(18)=>data_im_out(588),
            data_im_out(19)=>data_im_out(620),
            data_im_out(20)=>data_im_out(652),
            data_im_out(21)=>data_im_out(684),
            data_im_out(22)=>data_im_out(716),
            data_im_out(23)=>data_im_out(748),
            data_im_out(24)=>data_im_out(780),
            data_im_out(25)=>data_im_out(812),
            data_im_out(26)=>data_im_out(844),
            data_im_out(27)=>data_im_out(876),
            data_im_out(28)=>data_im_out(908),
            data_im_out(29)=>data_im_out(940),
            data_im_out(30)=>data_im_out(972),
            data_im_out(31)=>data_im_out(1004),
            data_im_out(32)=>data_im_out(1036),
            data_im_out(33)=>data_im_out(1068),
            data_im_out(34)=>data_im_out(1100),
            data_im_out(35)=>data_im_out(1132),
            data_im_out(36)=>data_im_out(1164),
            data_im_out(37)=>data_im_out(1196),
            data_im_out(38)=>data_im_out(1228),
            data_im_out(39)=>data_im_out(1260),
            data_im_out(40)=>data_im_out(1292),
            data_im_out(41)=>data_im_out(1324),
            data_im_out(42)=>data_im_out(1356),
            data_im_out(43)=>data_im_out(1388),
            data_im_out(44)=>data_im_out(1420),
            data_im_out(45)=>data_im_out(1452),
            data_im_out(46)=>data_im_out(1484),
            data_im_out(47)=>data_im_out(1516),
            data_im_out(48)=>data_im_out(1548),
            data_im_out(49)=>data_im_out(1580),
            data_im_out(50)=>data_im_out(1612),
            data_im_out(51)=>data_im_out(1644),
            data_im_out(52)=>data_im_out(1676),
            data_im_out(53)=>data_im_out(1708),
            data_im_out(54)=>data_im_out(1740),
            data_im_out(55)=>data_im_out(1772),
            data_im_out(56)=>data_im_out(1804),
            data_im_out(57)=>data_im_out(1836),
            data_im_out(58)=>data_im_out(1868),
            data_im_out(59)=>data_im_out(1900),
            data_im_out(60)=>data_im_out(1932),
            data_im_out(61)=>data_im_out(1964),
            data_im_out(62)=>data_im_out(1996),
            data_im_out(63)=>data_im_out(2028)
        );           

    URFFT_PT64_13 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(13),
            data_re_in(1)=>mul_re_out(45),
            data_re_in(2)=>mul_re_out(77),
            data_re_in(3)=>mul_re_out(109),
            data_re_in(4)=>mul_re_out(141),
            data_re_in(5)=>mul_re_out(173),
            data_re_in(6)=>mul_re_out(205),
            data_re_in(7)=>mul_re_out(237),
            data_re_in(8)=>mul_re_out(269),
            data_re_in(9)=>mul_re_out(301),
            data_re_in(10)=>mul_re_out(333),
            data_re_in(11)=>mul_re_out(365),
            data_re_in(12)=>mul_re_out(397),
            data_re_in(13)=>mul_re_out(429),
            data_re_in(14)=>mul_re_out(461),
            data_re_in(15)=>mul_re_out(493),
            data_re_in(16)=>mul_re_out(525),
            data_re_in(17)=>mul_re_out(557),
            data_re_in(18)=>mul_re_out(589),
            data_re_in(19)=>mul_re_out(621),
            data_re_in(20)=>mul_re_out(653),
            data_re_in(21)=>mul_re_out(685),
            data_re_in(22)=>mul_re_out(717),
            data_re_in(23)=>mul_re_out(749),
            data_re_in(24)=>mul_re_out(781),
            data_re_in(25)=>mul_re_out(813),
            data_re_in(26)=>mul_re_out(845),
            data_re_in(27)=>mul_re_out(877),
            data_re_in(28)=>mul_re_out(909),
            data_re_in(29)=>mul_re_out(941),
            data_re_in(30)=>mul_re_out(973),
            data_re_in(31)=>mul_re_out(1005),
            data_re_in(32)=>mul_re_out(1037),
            data_re_in(33)=>mul_re_out(1069),
            data_re_in(34)=>mul_re_out(1101),
            data_re_in(35)=>mul_re_out(1133),
            data_re_in(36)=>mul_re_out(1165),
            data_re_in(37)=>mul_re_out(1197),
            data_re_in(38)=>mul_re_out(1229),
            data_re_in(39)=>mul_re_out(1261),
            data_re_in(40)=>mul_re_out(1293),
            data_re_in(41)=>mul_re_out(1325),
            data_re_in(42)=>mul_re_out(1357),
            data_re_in(43)=>mul_re_out(1389),
            data_re_in(44)=>mul_re_out(1421),
            data_re_in(45)=>mul_re_out(1453),
            data_re_in(46)=>mul_re_out(1485),
            data_re_in(47)=>mul_re_out(1517),
            data_re_in(48)=>mul_re_out(1549),
            data_re_in(49)=>mul_re_out(1581),
            data_re_in(50)=>mul_re_out(1613),
            data_re_in(51)=>mul_re_out(1645),
            data_re_in(52)=>mul_re_out(1677),
            data_re_in(53)=>mul_re_out(1709),
            data_re_in(54)=>mul_re_out(1741),
            data_re_in(55)=>mul_re_out(1773),
            data_re_in(56)=>mul_re_out(1805),
            data_re_in(57)=>mul_re_out(1837),
            data_re_in(58)=>mul_re_out(1869),
            data_re_in(59)=>mul_re_out(1901),
            data_re_in(60)=>mul_re_out(1933),
            data_re_in(61)=>mul_re_out(1965),
            data_re_in(62)=>mul_re_out(1997),
            data_re_in(63)=>mul_re_out(2029),
            data_im_in(0)=>mul_im_out(13),
            data_im_in(1)=>mul_im_out(45),
            data_im_in(2)=>mul_im_out(77),
            data_im_in(3)=>mul_im_out(109),
            data_im_in(4)=>mul_im_out(141),
            data_im_in(5)=>mul_im_out(173),
            data_im_in(6)=>mul_im_out(205),
            data_im_in(7)=>mul_im_out(237),
            data_im_in(8)=>mul_im_out(269),
            data_im_in(9)=>mul_im_out(301),
            data_im_in(10)=>mul_im_out(333),
            data_im_in(11)=>mul_im_out(365),
            data_im_in(12)=>mul_im_out(397),
            data_im_in(13)=>mul_im_out(429),
            data_im_in(14)=>mul_im_out(461),
            data_im_in(15)=>mul_im_out(493),
            data_im_in(16)=>mul_im_out(525),
            data_im_in(17)=>mul_im_out(557),
            data_im_in(18)=>mul_im_out(589),
            data_im_in(19)=>mul_im_out(621),
            data_im_in(20)=>mul_im_out(653),
            data_im_in(21)=>mul_im_out(685),
            data_im_in(22)=>mul_im_out(717),
            data_im_in(23)=>mul_im_out(749),
            data_im_in(24)=>mul_im_out(781),
            data_im_in(25)=>mul_im_out(813),
            data_im_in(26)=>mul_im_out(845),
            data_im_in(27)=>mul_im_out(877),
            data_im_in(28)=>mul_im_out(909),
            data_im_in(29)=>mul_im_out(941),
            data_im_in(30)=>mul_im_out(973),
            data_im_in(31)=>mul_im_out(1005),
            data_im_in(32)=>mul_im_out(1037),
            data_im_in(33)=>mul_im_out(1069),
            data_im_in(34)=>mul_im_out(1101),
            data_im_in(35)=>mul_im_out(1133),
            data_im_in(36)=>mul_im_out(1165),
            data_im_in(37)=>mul_im_out(1197),
            data_im_in(38)=>mul_im_out(1229),
            data_im_in(39)=>mul_im_out(1261),
            data_im_in(40)=>mul_im_out(1293),
            data_im_in(41)=>mul_im_out(1325),
            data_im_in(42)=>mul_im_out(1357),
            data_im_in(43)=>mul_im_out(1389),
            data_im_in(44)=>mul_im_out(1421),
            data_im_in(45)=>mul_im_out(1453),
            data_im_in(46)=>mul_im_out(1485),
            data_im_in(47)=>mul_im_out(1517),
            data_im_in(48)=>mul_im_out(1549),
            data_im_in(49)=>mul_im_out(1581),
            data_im_in(50)=>mul_im_out(1613),
            data_im_in(51)=>mul_im_out(1645),
            data_im_in(52)=>mul_im_out(1677),
            data_im_in(53)=>mul_im_out(1709),
            data_im_in(54)=>mul_im_out(1741),
            data_im_in(55)=>mul_im_out(1773),
            data_im_in(56)=>mul_im_out(1805),
            data_im_in(57)=>mul_im_out(1837),
            data_im_in(58)=>mul_im_out(1869),
            data_im_in(59)=>mul_im_out(1901),
            data_im_in(60)=>mul_im_out(1933),
            data_im_in(61)=>mul_im_out(1965),
            data_im_in(62)=>mul_im_out(1997),
            data_im_in(63)=>mul_im_out(2029),
            data_re_out(0)=>data_re_out(13),
            data_re_out(1)=>data_re_out(45),
            data_re_out(2)=>data_re_out(77),
            data_re_out(3)=>data_re_out(109),
            data_re_out(4)=>data_re_out(141),
            data_re_out(5)=>data_re_out(173),
            data_re_out(6)=>data_re_out(205),
            data_re_out(7)=>data_re_out(237),
            data_re_out(8)=>data_re_out(269),
            data_re_out(9)=>data_re_out(301),
            data_re_out(10)=>data_re_out(333),
            data_re_out(11)=>data_re_out(365),
            data_re_out(12)=>data_re_out(397),
            data_re_out(13)=>data_re_out(429),
            data_re_out(14)=>data_re_out(461),
            data_re_out(15)=>data_re_out(493),
            data_re_out(16)=>data_re_out(525),
            data_re_out(17)=>data_re_out(557),
            data_re_out(18)=>data_re_out(589),
            data_re_out(19)=>data_re_out(621),
            data_re_out(20)=>data_re_out(653),
            data_re_out(21)=>data_re_out(685),
            data_re_out(22)=>data_re_out(717),
            data_re_out(23)=>data_re_out(749),
            data_re_out(24)=>data_re_out(781),
            data_re_out(25)=>data_re_out(813),
            data_re_out(26)=>data_re_out(845),
            data_re_out(27)=>data_re_out(877),
            data_re_out(28)=>data_re_out(909),
            data_re_out(29)=>data_re_out(941),
            data_re_out(30)=>data_re_out(973),
            data_re_out(31)=>data_re_out(1005),
            data_re_out(32)=>data_re_out(1037),
            data_re_out(33)=>data_re_out(1069),
            data_re_out(34)=>data_re_out(1101),
            data_re_out(35)=>data_re_out(1133),
            data_re_out(36)=>data_re_out(1165),
            data_re_out(37)=>data_re_out(1197),
            data_re_out(38)=>data_re_out(1229),
            data_re_out(39)=>data_re_out(1261),
            data_re_out(40)=>data_re_out(1293),
            data_re_out(41)=>data_re_out(1325),
            data_re_out(42)=>data_re_out(1357),
            data_re_out(43)=>data_re_out(1389),
            data_re_out(44)=>data_re_out(1421),
            data_re_out(45)=>data_re_out(1453),
            data_re_out(46)=>data_re_out(1485),
            data_re_out(47)=>data_re_out(1517),
            data_re_out(48)=>data_re_out(1549),
            data_re_out(49)=>data_re_out(1581),
            data_re_out(50)=>data_re_out(1613),
            data_re_out(51)=>data_re_out(1645),
            data_re_out(52)=>data_re_out(1677),
            data_re_out(53)=>data_re_out(1709),
            data_re_out(54)=>data_re_out(1741),
            data_re_out(55)=>data_re_out(1773),
            data_re_out(56)=>data_re_out(1805),
            data_re_out(57)=>data_re_out(1837),
            data_re_out(58)=>data_re_out(1869),
            data_re_out(59)=>data_re_out(1901),
            data_re_out(60)=>data_re_out(1933),
            data_re_out(61)=>data_re_out(1965),
            data_re_out(62)=>data_re_out(1997),
            data_re_out(63)=>data_re_out(2029),
            data_im_out(0)=>data_im_out(13),
            data_im_out(1)=>data_im_out(45),
            data_im_out(2)=>data_im_out(77),
            data_im_out(3)=>data_im_out(109),
            data_im_out(4)=>data_im_out(141),
            data_im_out(5)=>data_im_out(173),
            data_im_out(6)=>data_im_out(205),
            data_im_out(7)=>data_im_out(237),
            data_im_out(8)=>data_im_out(269),
            data_im_out(9)=>data_im_out(301),
            data_im_out(10)=>data_im_out(333),
            data_im_out(11)=>data_im_out(365),
            data_im_out(12)=>data_im_out(397),
            data_im_out(13)=>data_im_out(429),
            data_im_out(14)=>data_im_out(461),
            data_im_out(15)=>data_im_out(493),
            data_im_out(16)=>data_im_out(525),
            data_im_out(17)=>data_im_out(557),
            data_im_out(18)=>data_im_out(589),
            data_im_out(19)=>data_im_out(621),
            data_im_out(20)=>data_im_out(653),
            data_im_out(21)=>data_im_out(685),
            data_im_out(22)=>data_im_out(717),
            data_im_out(23)=>data_im_out(749),
            data_im_out(24)=>data_im_out(781),
            data_im_out(25)=>data_im_out(813),
            data_im_out(26)=>data_im_out(845),
            data_im_out(27)=>data_im_out(877),
            data_im_out(28)=>data_im_out(909),
            data_im_out(29)=>data_im_out(941),
            data_im_out(30)=>data_im_out(973),
            data_im_out(31)=>data_im_out(1005),
            data_im_out(32)=>data_im_out(1037),
            data_im_out(33)=>data_im_out(1069),
            data_im_out(34)=>data_im_out(1101),
            data_im_out(35)=>data_im_out(1133),
            data_im_out(36)=>data_im_out(1165),
            data_im_out(37)=>data_im_out(1197),
            data_im_out(38)=>data_im_out(1229),
            data_im_out(39)=>data_im_out(1261),
            data_im_out(40)=>data_im_out(1293),
            data_im_out(41)=>data_im_out(1325),
            data_im_out(42)=>data_im_out(1357),
            data_im_out(43)=>data_im_out(1389),
            data_im_out(44)=>data_im_out(1421),
            data_im_out(45)=>data_im_out(1453),
            data_im_out(46)=>data_im_out(1485),
            data_im_out(47)=>data_im_out(1517),
            data_im_out(48)=>data_im_out(1549),
            data_im_out(49)=>data_im_out(1581),
            data_im_out(50)=>data_im_out(1613),
            data_im_out(51)=>data_im_out(1645),
            data_im_out(52)=>data_im_out(1677),
            data_im_out(53)=>data_im_out(1709),
            data_im_out(54)=>data_im_out(1741),
            data_im_out(55)=>data_im_out(1773),
            data_im_out(56)=>data_im_out(1805),
            data_im_out(57)=>data_im_out(1837),
            data_im_out(58)=>data_im_out(1869),
            data_im_out(59)=>data_im_out(1901),
            data_im_out(60)=>data_im_out(1933),
            data_im_out(61)=>data_im_out(1965),
            data_im_out(62)=>data_im_out(1997),
            data_im_out(63)=>data_im_out(2029)
        );           

    URFFT_PT64_14 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(14),
            data_re_in(1)=>mul_re_out(46),
            data_re_in(2)=>mul_re_out(78),
            data_re_in(3)=>mul_re_out(110),
            data_re_in(4)=>mul_re_out(142),
            data_re_in(5)=>mul_re_out(174),
            data_re_in(6)=>mul_re_out(206),
            data_re_in(7)=>mul_re_out(238),
            data_re_in(8)=>mul_re_out(270),
            data_re_in(9)=>mul_re_out(302),
            data_re_in(10)=>mul_re_out(334),
            data_re_in(11)=>mul_re_out(366),
            data_re_in(12)=>mul_re_out(398),
            data_re_in(13)=>mul_re_out(430),
            data_re_in(14)=>mul_re_out(462),
            data_re_in(15)=>mul_re_out(494),
            data_re_in(16)=>mul_re_out(526),
            data_re_in(17)=>mul_re_out(558),
            data_re_in(18)=>mul_re_out(590),
            data_re_in(19)=>mul_re_out(622),
            data_re_in(20)=>mul_re_out(654),
            data_re_in(21)=>mul_re_out(686),
            data_re_in(22)=>mul_re_out(718),
            data_re_in(23)=>mul_re_out(750),
            data_re_in(24)=>mul_re_out(782),
            data_re_in(25)=>mul_re_out(814),
            data_re_in(26)=>mul_re_out(846),
            data_re_in(27)=>mul_re_out(878),
            data_re_in(28)=>mul_re_out(910),
            data_re_in(29)=>mul_re_out(942),
            data_re_in(30)=>mul_re_out(974),
            data_re_in(31)=>mul_re_out(1006),
            data_re_in(32)=>mul_re_out(1038),
            data_re_in(33)=>mul_re_out(1070),
            data_re_in(34)=>mul_re_out(1102),
            data_re_in(35)=>mul_re_out(1134),
            data_re_in(36)=>mul_re_out(1166),
            data_re_in(37)=>mul_re_out(1198),
            data_re_in(38)=>mul_re_out(1230),
            data_re_in(39)=>mul_re_out(1262),
            data_re_in(40)=>mul_re_out(1294),
            data_re_in(41)=>mul_re_out(1326),
            data_re_in(42)=>mul_re_out(1358),
            data_re_in(43)=>mul_re_out(1390),
            data_re_in(44)=>mul_re_out(1422),
            data_re_in(45)=>mul_re_out(1454),
            data_re_in(46)=>mul_re_out(1486),
            data_re_in(47)=>mul_re_out(1518),
            data_re_in(48)=>mul_re_out(1550),
            data_re_in(49)=>mul_re_out(1582),
            data_re_in(50)=>mul_re_out(1614),
            data_re_in(51)=>mul_re_out(1646),
            data_re_in(52)=>mul_re_out(1678),
            data_re_in(53)=>mul_re_out(1710),
            data_re_in(54)=>mul_re_out(1742),
            data_re_in(55)=>mul_re_out(1774),
            data_re_in(56)=>mul_re_out(1806),
            data_re_in(57)=>mul_re_out(1838),
            data_re_in(58)=>mul_re_out(1870),
            data_re_in(59)=>mul_re_out(1902),
            data_re_in(60)=>mul_re_out(1934),
            data_re_in(61)=>mul_re_out(1966),
            data_re_in(62)=>mul_re_out(1998),
            data_re_in(63)=>mul_re_out(2030),
            data_im_in(0)=>mul_im_out(14),
            data_im_in(1)=>mul_im_out(46),
            data_im_in(2)=>mul_im_out(78),
            data_im_in(3)=>mul_im_out(110),
            data_im_in(4)=>mul_im_out(142),
            data_im_in(5)=>mul_im_out(174),
            data_im_in(6)=>mul_im_out(206),
            data_im_in(7)=>mul_im_out(238),
            data_im_in(8)=>mul_im_out(270),
            data_im_in(9)=>mul_im_out(302),
            data_im_in(10)=>mul_im_out(334),
            data_im_in(11)=>mul_im_out(366),
            data_im_in(12)=>mul_im_out(398),
            data_im_in(13)=>mul_im_out(430),
            data_im_in(14)=>mul_im_out(462),
            data_im_in(15)=>mul_im_out(494),
            data_im_in(16)=>mul_im_out(526),
            data_im_in(17)=>mul_im_out(558),
            data_im_in(18)=>mul_im_out(590),
            data_im_in(19)=>mul_im_out(622),
            data_im_in(20)=>mul_im_out(654),
            data_im_in(21)=>mul_im_out(686),
            data_im_in(22)=>mul_im_out(718),
            data_im_in(23)=>mul_im_out(750),
            data_im_in(24)=>mul_im_out(782),
            data_im_in(25)=>mul_im_out(814),
            data_im_in(26)=>mul_im_out(846),
            data_im_in(27)=>mul_im_out(878),
            data_im_in(28)=>mul_im_out(910),
            data_im_in(29)=>mul_im_out(942),
            data_im_in(30)=>mul_im_out(974),
            data_im_in(31)=>mul_im_out(1006),
            data_im_in(32)=>mul_im_out(1038),
            data_im_in(33)=>mul_im_out(1070),
            data_im_in(34)=>mul_im_out(1102),
            data_im_in(35)=>mul_im_out(1134),
            data_im_in(36)=>mul_im_out(1166),
            data_im_in(37)=>mul_im_out(1198),
            data_im_in(38)=>mul_im_out(1230),
            data_im_in(39)=>mul_im_out(1262),
            data_im_in(40)=>mul_im_out(1294),
            data_im_in(41)=>mul_im_out(1326),
            data_im_in(42)=>mul_im_out(1358),
            data_im_in(43)=>mul_im_out(1390),
            data_im_in(44)=>mul_im_out(1422),
            data_im_in(45)=>mul_im_out(1454),
            data_im_in(46)=>mul_im_out(1486),
            data_im_in(47)=>mul_im_out(1518),
            data_im_in(48)=>mul_im_out(1550),
            data_im_in(49)=>mul_im_out(1582),
            data_im_in(50)=>mul_im_out(1614),
            data_im_in(51)=>mul_im_out(1646),
            data_im_in(52)=>mul_im_out(1678),
            data_im_in(53)=>mul_im_out(1710),
            data_im_in(54)=>mul_im_out(1742),
            data_im_in(55)=>mul_im_out(1774),
            data_im_in(56)=>mul_im_out(1806),
            data_im_in(57)=>mul_im_out(1838),
            data_im_in(58)=>mul_im_out(1870),
            data_im_in(59)=>mul_im_out(1902),
            data_im_in(60)=>mul_im_out(1934),
            data_im_in(61)=>mul_im_out(1966),
            data_im_in(62)=>mul_im_out(1998),
            data_im_in(63)=>mul_im_out(2030),
            data_re_out(0)=>data_re_out(14),
            data_re_out(1)=>data_re_out(46),
            data_re_out(2)=>data_re_out(78),
            data_re_out(3)=>data_re_out(110),
            data_re_out(4)=>data_re_out(142),
            data_re_out(5)=>data_re_out(174),
            data_re_out(6)=>data_re_out(206),
            data_re_out(7)=>data_re_out(238),
            data_re_out(8)=>data_re_out(270),
            data_re_out(9)=>data_re_out(302),
            data_re_out(10)=>data_re_out(334),
            data_re_out(11)=>data_re_out(366),
            data_re_out(12)=>data_re_out(398),
            data_re_out(13)=>data_re_out(430),
            data_re_out(14)=>data_re_out(462),
            data_re_out(15)=>data_re_out(494),
            data_re_out(16)=>data_re_out(526),
            data_re_out(17)=>data_re_out(558),
            data_re_out(18)=>data_re_out(590),
            data_re_out(19)=>data_re_out(622),
            data_re_out(20)=>data_re_out(654),
            data_re_out(21)=>data_re_out(686),
            data_re_out(22)=>data_re_out(718),
            data_re_out(23)=>data_re_out(750),
            data_re_out(24)=>data_re_out(782),
            data_re_out(25)=>data_re_out(814),
            data_re_out(26)=>data_re_out(846),
            data_re_out(27)=>data_re_out(878),
            data_re_out(28)=>data_re_out(910),
            data_re_out(29)=>data_re_out(942),
            data_re_out(30)=>data_re_out(974),
            data_re_out(31)=>data_re_out(1006),
            data_re_out(32)=>data_re_out(1038),
            data_re_out(33)=>data_re_out(1070),
            data_re_out(34)=>data_re_out(1102),
            data_re_out(35)=>data_re_out(1134),
            data_re_out(36)=>data_re_out(1166),
            data_re_out(37)=>data_re_out(1198),
            data_re_out(38)=>data_re_out(1230),
            data_re_out(39)=>data_re_out(1262),
            data_re_out(40)=>data_re_out(1294),
            data_re_out(41)=>data_re_out(1326),
            data_re_out(42)=>data_re_out(1358),
            data_re_out(43)=>data_re_out(1390),
            data_re_out(44)=>data_re_out(1422),
            data_re_out(45)=>data_re_out(1454),
            data_re_out(46)=>data_re_out(1486),
            data_re_out(47)=>data_re_out(1518),
            data_re_out(48)=>data_re_out(1550),
            data_re_out(49)=>data_re_out(1582),
            data_re_out(50)=>data_re_out(1614),
            data_re_out(51)=>data_re_out(1646),
            data_re_out(52)=>data_re_out(1678),
            data_re_out(53)=>data_re_out(1710),
            data_re_out(54)=>data_re_out(1742),
            data_re_out(55)=>data_re_out(1774),
            data_re_out(56)=>data_re_out(1806),
            data_re_out(57)=>data_re_out(1838),
            data_re_out(58)=>data_re_out(1870),
            data_re_out(59)=>data_re_out(1902),
            data_re_out(60)=>data_re_out(1934),
            data_re_out(61)=>data_re_out(1966),
            data_re_out(62)=>data_re_out(1998),
            data_re_out(63)=>data_re_out(2030),
            data_im_out(0)=>data_im_out(14),
            data_im_out(1)=>data_im_out(46),
            data_im_out(2)=>data_im_out(78),
            data_im_out(3)=>data_im_out(110),
            data_im_out(4)=>data_im_out(142),
            data_im_out(5)=>data_im_out(174),
            data_im_out(6)=>data_im_out(206),
            data_im_out(7)=>data_im_out(238),
            data_im_out(8)=>data_im_out(270),
            data_im_out(9)=>data_im_out(302),
            data_im_out(10)=>data_im_out(334),
            data_im_out(11)=>data_im_out(366),
            data_im_out(12)=>data_im_out(398),
            data_im_out(13)=>data_im_out(430),
            data_im_out(14)=>data_im_out(462),
            data_im_out(15)=>data_im_out(494),
            data_im_out(16)=>data_im_out(526),
            data_im_out(17)=>data_im_out(558),
            data_im_out(18)=>data_im_out(590),
            data_im_out(19)=>data_im_out(622),
            data_im_out(20)=>data_im_out(654),
            data_im_out(21)=>data_im_out(686),
            data_im_out(22)=>data_im_out(718),
            data_im_out(23)=>data_im_out(750),
            data_im_out(24)=>data_im_out(782),
            data_im_out(25)=>data_im_out(814),
            data_im_out(26)=>data_im_out(846),
            data_im_out(27)=>data_im_out(878),
            data_im_out(28)=>data_im_out(910),
            data_im_out(29)=>data_im_out(942),
            data_im_out(30)=>data_im_out(974),
            data_im_out(31)=>data_im_out(1006),
            data_im_out(32)=>data_im_out(1038),
            data_im_out(33)=>data_im_out(1070),
            data_im_out(34)=>data_im_out(1102),
            data_im_out(35)=>data_im_out(1134),
            data_im_out(36)=>data_im_out(1166),
            data_im_out(37)=>data_im_out(1198),
            data_im_out(38)=>data_im_out(1230),
            data_im_out(39)=>data_im_out(1262),
            data_im_out(40)=>data_im_out(1294),
            data_im_out(41)=>data_im_out(1326),
            data_im_out(42)=>data_im_out(1358),
            data_im_out(43)=>data_im_out(1390),
            data_im_out(44)=>data_im_out(1422),
            data_im_out(45)=>data_im_out(1454),
            data_im_out(46)=>data_im_out(1486),
            data_im_out(47)=>data_im_out(1518),
            data_im_out(48)=>data_im_out(1550),
            data_im_out(49)=>data_im_out(1582),
            data_im_out(50)=>data_im_out(1614),
            data_im_out(51)=>data_im_out(1646),
            data_im_out(52)=>data_im_out(1678),
            data_im_out(53)=>data_im_out(1710),
            data_im_out(54)=>data_im_out(1742),
            data_im_out(55)=>data_im_out(1774),
            data_im_out(56)=>data_im_out(1806),
            data_im_out(57)=>data_im_out(1838),
            data_im_out(58)=>data_im_out(1870),
            data_im_out(59)=>data_im_out(1902),
            data_im_out(60)=>data_im_out(1934),
            data_im_out(61)=>data_im_out(1966),
            data_im_out(62)=>data_im_out(1998),
            data_im_out(63)=>data_im_out(2030)
        );           

    URFFT_PT64_15 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(15),
            data_re_in(1)=>mul_re_out(47),
            data_re_in(2)=>mul_re_out(79),
            data_re_in(3)=>mul_re_out(111),
            data_re_in(4)=>mul_re_out(143),
            data_re_in(5)=>mul_re_out(175),
            data_re_in(6)=>mul_re_out(207),
            data_re_in(7)=>mul_re_out(239),
            data_re_in(8)=>mul_re_out(271),
            data_re_in(9)=>mul_re_out(303),
            data_re_in(10)=>mul_re_out(335),
            data_re_in(11)=>mul_re_out(367),
            data_re_in(12)=>mul_re_out(399),
            data_re_in(13)=>mul_re_out(431),
            data_re_in(14)=>mul_re_out(463),
            data_re_in(15)=>mul_re_out(495),
            data_re_in(16)=>mul_re_out(527),
            data_re_in(17)=>mul_re_out(559),
            data_re_in(18)=>mul_re_out(591),
            data_re_in(19)=>mul_re_out(623),
            data_re_in(20)=>mul_re_out(655),
            data_re_in(21)=>mul_re_out(687),
            data_re_in(22)=>mul_re_out(719),
            data_re_in(23)=>mul_re_out(751),
            data_re_in(24)=>mul_re_out(783),
            data_re_in(25)=>mul_re_out(815),
            data_re_in(26)=>mul_re_out(847),
            data_re_in(27)=>mul_re_out(879),
            data_re_in(28)=>mul_re_out(911),
            data_re_in(29)=>mul_re_out(943),
            data_re_in(30)=>mul_re_out(975),
            data_re_in(31)=>mul_re_out(1007),
            data_re_in(32)=>mul_re_out(1039),
            data_re_in(33)=>mul_re_out(1071),
            data_re_in(34)=>mul_re_out(1103),
            data_re_in(35)=>mul_re_out(1135),
            data_re_in(36)=>mul_re_out(1167),
            data_re_in(37)=>mul_re_out(1199),
            data_re_in(38)=>mul_re_out(1231),
            data_re_in(39)=>mul_re_out(1263),
            data_re_in(40)=>mul_re_out(1295),
            data_re_in(41)=>mul_re_out(1327),
            data_re_in(42)=>mul_re_out(1359),
            data_re_in(43)=>mul_re_out(1391),
            data_re_in(44)=>mul_re_out(1423),
            data_re_in(45)=>mul_re_out(1455),
            data_re_in(46)=>mul_re_out(1487),
            data_re_in(47)=>mul_re_out(1519),
            data_re_in(48)=>mul_re_out(1551),
            data_re_in(49)=>mul_re_out(1583),
            data_re_in(50)=>mul_re_out(1615),
            data_re_in(51)=>mul_re_out(1647),
            data_re_in(52)=>mul_re_out(1679),
            data_re_in(53)=>mul_re_out(1711),
            data_re_in(54)=>mul_re_out(1743),
            data_re_in(55)=>mul_re_out(1775),
            data_re_in(56)=>mul_re_out(1807),
            data_re_in(57)=>mul_re_out(1839),
            data_re_in(58)=>mul_re_out(1871),
            data_re_in(59)=>mul_re_out(1903),
            data_re_in(60)=>mul_re_out(1935),
            data_re_in(61)=>mul_re_out(1967),
            data_re_in(62)=>mul_re_out(1999),
            data_re_in(63)=>mul_re_out(2031),
            data_im_in(0)=>mul_im_out(15),
            data_im_in(1)=>mul_im_out(47),
            data_im_in(2)=>mul_im_out(79),
            data_im_in(3)=>mul_im_out(111),
            data_im_in(4)=>mul_im_out(143),
            data_im_in(5)=>mul_im_out(175),
            data_im_in(6)=>mul_im_out(207),
            data_im_in(7)=>mul_im_out(239),
            data_im_in(8)=>mul_im_out(271),
            data_im_in(9)=>mul_im_out(303),
            data_im_in(10)=>mul_im_out(335),
            data_im_in(11)=>mul_im_out(367),
            data_im_in(12)=>mul_im_out(399),
            data_im_in(13)=>mul_im_out(431),
            data_im_in(14)=>mul_im_out(463),
            data_im_in(15)=>mul_im_out(495),
            data_im_in(16)=>mul_im_out(527),
            data_im_in(17)=>mul_im_out(559),
            data_im_in(18)=>mul_im_out(591),
            data_im_in(19)=>mul_im_out(623),
            data_im_in(20)=>mul_im_out(655),
            data_im_in(21)=>mul_im_out(687),
            data_im_in(22)=>mul_im_out(719),
            data_im_in(23)=>mul_im_out(751),
            data_im_in(24)=>mul_im_out(783),
            data_im_in(25)=>mul_im_out(815),
            data_im_in(26)=>mul_im_out(847),
            data_im_in(27)=>mul_im_out(879),
            data_im_in(28)=>mul_im_out(911),
            data_im_in(29)=>mul_im_out(943),
            data_im_in(30)=>mul_im_out(975),
            data_im_in(31)=>mul_im_out(1007),
            data_im_in(32)=>mul_im_out(1039),
            data_im_in(33)=>mul_im_out(1071),
            data_im_in(34)=>mul_im_out(1103),
            data_im_in(35)=>mul_im_out(1135),
            data_im_in(36)=>mul_im_out(1167),
            data_im_in(37)=>mul_im_out(1199),
            data_im_in(38)=>mul_im_out(1231),
            data_im_in(39)=>mul_im_out(1263),
            data_im_in(40)=>mul_im_out(1295),
            data_im_in(41)=>mul_im_out(1327),
            data_im_in(42)=>mul_im_out(1359),
            data_im_in(43)=>mul_im_out(1391),
            data_im_in(44)=>mul_im_out(1423),
            data_im_in(45)=>mul_im_out(1455),
            data_im_in(46)=>mul_im_out(1487),
            data_im_in(47)=>mul_im_out(1519),
            data_im_in(48)=>mul_im_out(1551),
            data_im_in(49)=>mul_im_out(1583),
            data_im_in(50)=>mul_im_out(1615),
            data_im_in(51)=>mul_im_out(1647),
            data_im_in(52)=>mul_im_out(1679),
            data_im_in(53)=>mul_im_out(1711),
            data_im_in(54)=>mul_im_out(1743),
            data_im_in(55)=>mul_im_out(1775),
            data_im_in(56)=>mul_im_out(1807),
            data_im_in(57)=>mul_im_out(1839),
            data_im_in(58)=>mul_im_out(1871),
            data_im_in(59)=>mul_im_out(1903),
            data_im_in(60)=>mul_im_out(1935),
            data_im_in(61)=>mul_im_out(1967),
            data_im_in(62)=>mul_im_out(1999),
            data_im_in(63)=>mul_im_out(2031),
            data_re_out(0)=>data_re_out(15),
            data_re_out(1)=>data_re_out(47),
            data_re_out(2)=>data_re_out(79),
            data_re_out(3)=>data_re_out(111),
            data_re_out(4)=>data_re_out(143),
            data_re_out(5)=>data_re_out(175),
            data_re_out(6)=>data_re_out(207),
            data_re_out(7)=>data_re_out(239),
            data_re_out(8)=>data_re_out(271),
            data_re_out(9)=>data_re_out(303),
            data_re_out(10)=>data_re_out(335),
            data_re_out(11)=>data_re_out(367),
            data_re_out(12)=>data_re_out(399),
            data_re_out(13)=>data_re_out(431),
            data_re_out(14)=>data_re_out(463),
            data_re_out(15)=>data_re_out(495),
            data_re_out(16)=>data_re_out(527),
            data_re_out(17)=>data_re_out(559),
            data_re_out(18)=>data_re_out(591),
            data_re_out(19)=>data_re_out(623),
            data_re_out(20)=>data_re_out(655),
            data_re_out(21)=>data_re_out(687),
            data_re_out(22)=>data_re_out(719),
            data_re_out(23)=>data_re_out(751),
            data_re_out(24)=>data_re_out(783),
            data_re_out(25)=>data_re_out(815),
            data_re_out(26)=>data_re_out(847),
            data_re_out(27)=>data_re_out(879),
            data_re_out(28)=>data_re_out(911),
            data_re_out(29)=>data_re_out(943),
            data_re_out(30)=>data_re_out(975),
            data_re_out(31)=>data_re_out(1007),
            data_re_out(32)=>data_re_out(1039),
            data_re_out(33)=>data_re_out(1071),
            data_re_out(34)=>data_re_out(1103),
            data_re_out(35)=>data_re_out(1135),
            data_re_out(36)=>data_re_out(1167),
            data_re_out(37)=>data_re_out(1199),
            data_re_out(38)=>data_re_out(1231),
            data_re_out(39)=>data_re_out(1263),
            data_re_out(40)=>data_re_out(1295),
            data_re_out(41)=>data_re_out(1327),
            data_re_out(42)=>data_re_out(1359),
            data_re_out(43)=>data_re_out(1391),
            data_re_out(44)=>data_re_out(1423),
            data_re_out(45)=>data_re_out(1455),
            data_re_out(46)=>data_re_out(1487),
            data_re_out(47)=>data_re_out(1519),
            data_re_out(48)=>data_re_out(1551),
            data_re_out(49)=>data_re_out(1583),
            data_re_out(50)=>data_re_out(1615),
            data_re_out(51)=>data_re_out(1647),
            data_re_out(52)=>data_re_out(1679),
            data_re_out(53)=>data_re_out(1711),
            data_re_out(54)=>data_re_out(1743),
            data_re_out(55)=>data_re_out(1775),
            data_re_out(56)=>data_re_out(1807),
            data_re_out(57)=>data_re_out(1839),
            data_re_out(58)=>data_re_out(1871),
            data_re_out(59)=>data_re_out(1903),
            data_re_out(60)=>data_re_out(1935),
            data_re_out(61)=>data_re_out(1967),
            data_re_out(62)=>data_re_out(1999),
            data_re_out(63)=>data_re_out(2031),
            data_im_out(0)=>data_im_out(15),
            data_im_out(1)=>data_im_out(47),
            data_im_out(2)=>data_im_out(79),
            data_im_out(3)=>data_im_out(111),
            data_im_out(4)=>data_im_out(143),
            data_im_out(5)=>data_im_out(175),
            data_im_out(6)=>data_im_out(207),
            data_im_out(7)=>data_im_out(239),
            data_im_out(8)=>data_im_out(271),
            data_im_out(9)=>data_im_out(303),
            data_im_out(10)=>data_im_out(335),
            data_im_out(11)=>data_im_out(367),
            data_im_out(12)=>data_im_out(399),
            data_im_out(13)=>data_im_out(431),
            data_im_out(14)=>data_im_out(463),
            data_im_out(15)=>data_im_out(495),
            data_im_out(16)=>data_im_out(527),
            data_im_out(17)=>data_im_out(559),
            data_im_out(18)=>data_im_out(591),
            data_im_out(19)=>data_im_out(623),
            data_im_out(20)=>data_im_out(655),
            data_im_out(21)=>data_im_out(687),
            data_im_out(22)=>data_im_out(719),
            data_im_out(23)=>data_im_out(751),
            data_im_out(24)=>data_im_out(783),
            data_im_out(25)=>data_im_out(815),
            data_im_out(26)=>data_im_out(847),
            data_im_out(27)=>data_im_out(879),
            data_im_out(28)=>data_im_out(911),
            data_im_out(29)=>data_im_out(943),
            data_im_out(30)=>data_im_out(975),
            data_im_out(31)=>data_im_out(1007),
            data_im_out(32)=>data_im_out(1039),
            data_im_out(33)=>data_im_out(1071),
            data_im_out(34)=>data_im_out(1103),
            data_im_out(35)=>data_im_out(1135),
            data_im_out(36)=>data_im_out(1167),
            data_im_out(37)=>data_im_out(1199),
            data_im_out(38)=>data_im_out(1231),
            data_im_out(39)=>data_im_out(1263),
            data_im_out(40)=>data_im_out(1295),
            data_im_out(41)=>data_im_out(1327),
            data_im_out(42)=>data_im_out(1359),
            data_im_out(43)=>data_im_out(1391),
            data_im_out(44)=>data_im_out(1423),
            data_im_out(45)=>data_im_out(1455),
            data_im_out(46)=>data_im_out(1487),
            data_im_out(47)=>data_im_out(1519),
            data_im_out(48)=>data_im_out(1551),
            data_im_out(49)=>data_im_out(1583),
            data_im_out(50)=>data_im_out(1615),
            data_im_out(51)=>data_im_out(1647),
            data_im_out(52)=>data_im_out(1679),
            data_im_out(53)=>data_im_out(1711),
            data_im_out(54)=>data_im_out(1743),
            data_im_out(55)=>data_im_out(1775),
            data_im_out(56)=>data_im_out(1807),
            data_im_out(57)=>data_im_out(1839),
            data_im_out(58)=>data_im_out(1871),
            data_im_out(59)=>data_im_out(1903),
            data_im_out(60)=>data_im_out(1935),
            data_im_out(61)=>data_im_out(1967),
            data_im_out(62)=>data_im_out(1999),
            data_im_out(63)=>data_im_out(2031)
        );           

    URFFT_PT64_16 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(16),
            data_re_in(1)=>mul_re_out(48),
            data_re_in(2)=>mul_re_out(80),
            data_re_in(3)=>mul_re_out(112),
            data_re_in(4)=>mul_re_out(144),
            data_re_in(5)=>mul_re_out(176),
            data_re_in(6)=>mul_re_out(208),
            data_re_in(7)=>mul_re_out(240),
            data_re_in(8)=>mul_re_out(272),
            data_re_in(9)=>mul_re_out(304),
            data_re_in(10)=>mul_re_out(336),
            data_re_in(11)=>mul_re_out(368),
            data_re_in(12)=>mul_re_out(400),
            data_re_in(13)=>mul_re_out(432),
            data_re_in(14)=>mul_re_out(464),
            data_re_in(15)=>mul_re_out(496),
            data_re_in(16)=>mul_re_out(528),
            data_re_in(17)=>mul_re_out(560),
            data_re_in(18)=>mul_re_out(592),
            data_re_in(19)=>mul_re_out(624),
            data_re_in(20)=>mul_re_out(656),
            data_re_in(21)=>mul_re_out(688),
            data_re_in(22)=>mul_re_out(720),
            data_re_in(23)=>mul_re_out(752),
            data_re_in(24)=>mul_re_out(784),
            data_re_in(25)=>mul_re_out(816),
            data_re_in(26)=>mul_re_out(848),
            data_re_in(27)=>mul_re_out(880),
            data_re_in(28)=>mul_re_out(912),
            data_re_in(29)=>mul_re_out(944),
            data_re_in(30)=>mul_re_out(976),
            data_re_in(31)=>mul_re_out(1008),
            data_re_in(32)=>mul_re_out(1040),
            data_re_in(33)=>mul_re_out(1072),
            data_re_in(34)=>mul_re_out(1104),
            data_re_in(35)=>mul_re_out(1136),
            data_re_in(36)=>mul_re_out(1168),
            data_re_in(37)=>mul_re_out(1200),
            data_re_in(38)=>mul_re_out(1232),
            data_re_in(39)=>mul_re_out(1264),
            data_re_in(40)=>mul_re_out(1296),
            data_re_in(41)=>mul_re_out(1328),
            data_re_in(42)=>mul_re_out(1360),
            data_re_in(43)=>mul_re_out(1392),
            data_re_in(44)=>mul_re_out(1424),
            data_re_in(45)=>mul_re_out(1456),
            data_re_in(46)=>mul_re_out(1488),
            data_re_in(47)=>mul_re_out(1520),
            data_re_in(48)=>mul_re_out(1552),
            data_re_in(49)=>mul_re_out(1584),
            data_re_in(50)=>mul_re_out(1616),
            data_re_in(51)=>mul_re_out(1648),
            data_re_in(52)=>mul_re_out(1680),
            data_re_in(53)=>mul_re_out(1712),
            data_re_in(54)=>mul_re_out(1744),
            data_re_in(55)=>mul_re_out(1776),
            data_re_in(56)=>mul_re_out(1808),
            data_re_in(57)=>mul_re_out(1840),
            data_re_in(58)=>mul_re_out(1872),
            data_re_in(59)=>mul_re_out(1904),
            data_re_in(60)=>mul_re_out(1936),
            data_re_in(61)=>mul_re_out(1968),
            data_re_in(62)=>mul_re_out(2000),
            data_re_in(63)=>mul_re_out(2032),
            data_im_in(0)=>mul_im_out(16),
            data_im_in(1)=>mul_im_out(48),
            data_im_in(2)=>mul_im_out(80),
            data_im_in(3)=>mul_im_out(112),
            data_im_in(4)=>mul_im_out(144),
            data_im_in(5)=>mul_im_out(176),
            data_im_in(6)=>mul_im_out(208),
            data_im_in(7)=>mul_im_out(240),
            data_im_in(8)=>mul_im_out(272),
            data_im_in(9)=>mul_im_out(304),
            data_im_in(10)=>mul_im_out(336),
            data_im_in(11)=>mul_im_out(368),
            data_im_in(12)=>mul_im_out(400),
            data_im_in(13)=>mul_im_out(432),
            data_im_in(14)=>mul_im_out(464),
            data_im_in(15)=>mul_im_out(496),
            data_im_in(16)=>mul_im_out(528),
            data_im_in(17)=>mul_im_out(560),
            data_im_in(18)=>mul_im_out(592),
            data_im_in(19)=>mul_im_out(624),
            data_im_in(20)=>mul_im_out(656),
            data_im_in(21)=>mul_im_out(688),
            data_im_in(22)=>mul_im_out(720),
            data_im_in(23)=>mul_im_out(752),
            data_im_in(24)=>mul_im_out(784),
            data_im_in(25)=>mul_im_out(816),
            data_im_in(26)=>mul_im_out(848),
            data_im_in(27)=>mul_im_out(880),
            data_im_in(28)=>mul_im_out(912),
            data_im_in(29)=>mul_im_out(944),
            data_im_in(30)=>mul_im_out(976),
            data_im_in(31)=>mul_im_out(1008),
            data_im_in(32)=>mul_im_out(1040),
            data_im_in(33)=>mul_im_out(1072),
            data_im_in(34)=>mul_im_out(1104),
            data_im_in(35)=>mul_im_out(1136),
            data_im_in(36)=>mul_im_out(1168),
            data_im_in(37)=>mul_im_out(1200),
            data_im_in(38)=>mul_im_out(1232),
            data_im_in(39)=>mul_im_out(1264),
            data_im_in(40)=>mul_im_out(1296),
            data_im_in(41)=>mul_im_out(1328),
            data_im_in(42)=>mul_im_out(1360),
            data_im_in(43)=>mul_im_out(1392),
            data_im_in(44)=>mul_im_out(1424),
            data_im_in(45)=>mul_im_out(1456),
            data_im_in(46)=>mul_im_out(1488),
            data_im_in(47)=>mul_im_out(1520),
            data_im_in(48)=>mul_im_out(1552),
            data_im_in(49)=>mul_im_out(1584),
            data_im_in(50)=>mul_im_out(1616),
            data_im_in(51)=>mul_im_out(1648),
            data_im_in(52)=>mul_im_out(1680),
            data_im_in(53)=>mul_im_out(1712),
            data_im_in(54)=>mul_im_out(1744),
            data_im_in(55)=>mul_im_out(1776),
            data_im_in(56)=>mul_im_out(1808),
            data_im_in(57)=>mul_im_out(1840),
            data_im_in(58)=>mul_im_out(1872),
            data_im_in(59)=>mul_im_out(1904),
            data_im_in(60)=>mul_im_out(1936),
            data_im_in(61)=>mul_im_out(1968),
            data_im_in(62)=>mul_im_out(2000),
            data_im_in(63)=>mul_im_out(2032),
            data_re_out(0)=>data_re_out(16),
            data_re_out(1)=>data_re_out(48),
            data_re_out(2)=>data_re_out(80),
            data_re_out(3)=>data_re_out(112),
            data_re_out(4)=>data_re_out(144),
            data_re_out(5)=>data_re_out(176),
            data_re_out(6)=>data_re_out(208),
            data_re_out(7)=>data_re_out(240),
            data_re_out(8)=>data_re_out(272),
            data_re_out(9)=>data_re_out(304),
            data_re_out(10)=>data_re_out(336),
            data_re_out(11)=>data_re_out(368),
            data_re_out(12)=>data_re_out(400),
            data_re_out(13)=>data_re_out(432),
            data_re_out(14)=>data_re_out(464),
            data_re_out(15)=>data_re_out(496),
            data_re_out(16)=>data_re_out(528),
            data_re_out(17)=>data_re_out(560),
            data_re_out(18)=>data_re_out(592),
            data_re_out(19)=>data_re_out(624),
            data_re_out(20)=>data_re_out(656),
            data_re_out(21)=>data_re_out(688),
            data_re_out(22)=>data_re_out(720),
            data_re_out(23)=>data_re_out(752),
            data_re_out(24)=>data_re_out(784),
            data_re_out(25)=>data_re_out(816),
            data_re_out(26)=>data_re_out(848),
            data_re_out(27)=>data_re_out(880),
            data_re_out(28)=>data_re_out(912),
            data_re_out(29)=>data_re_out(944),
            data_re_out(30)=>data_re_out(976),
            data_re_out(31)=>data_re_out(1008),
            data_re_out(32)=>data_re_out(1040),
            data_re_out(33)=>data_re_out(1072),
            data_re_out(34)=>data_re_out(1104),
            data_re_out(35)=>data_re_out(1136),
            data_re_out(36)=>data_re_out(1168),
            data_re_out(37)=>data_re_out(1200),
            data_re_out(38)=>data_re_out(1232),
            data_re_out(39)=>data_re_out(1264),
            data_re_out(40)=>data_re_out(1296),
            data_re_out(41)=>data_re_out(1328),
            data_re_out(42)=>data_re_out(1360),
            data_re_out(43)=>data_re_out(1392),
            data_re_out(44)=>data_re_out(1424),
            data_re_out(45)=>data_re_out(1456),
            data_re_out(46)=>data_re_out(1488),
            data_re_out(47)=>data_re_out(1520),
            data_re_out(48)=>data_re_out(1552),
            data_re_out(49)=>data_re_out(1584),
            data_re_out(50)=>data_re_out(1616),
            data_re_out(51)=>data_re_out(1648),
            data_re_out(52)=>data_re_out(1680),
            data_re_out(53)=>data_re_out(1712),
            data_re_out(54)=>data_re_out(1744),
            data_re_out(55)=>data_re_out(1776),
            data_re_out(56)=>data_re_out(1808),
            data_re_out(57)=>data_re_out(1840),
            data_re_out(58)=>data_re_out(1872),
            data_re_out(59)=>data_re_out(1904),
            data_re_out(60)=>data_re_out(1936),
            data_re_out(61)=>data_re_out(1968),
            data_re_out(62)=>data_re_out(2000),
            data_re_out(63)=>data_re_out(2032),
            data_im_out(0)=>data_im_out(16),
            data_im_out(1)=>data_im_out(48),
            data_im_out(2)=>data_im_out(80),
            data_im_out(3)=>data_im_out(112),
            data_im_out(4)=>data_im_out(144),
            data_im_out(5)=>data_im_out(176),
            data_im_out(6)=>data_im_out(208),
            data_im_out(7)=>data_im_out(240),
            data_im_out(8)=>data_im_out(272),
            data_im_out(9)=>data_im_out(304),
            data_im_out(10)=>data_im_out(336),
            data_im_out(11)=>data_im_out(368),
            data_im_out(12)=>data_im_out(400),
            data_im_out(13)=>data_im_out(432),
            data_im_out(14)=>data_im_out(464),
            data_im_out(15)=>data_im_out(496),
            data_im_out(16)=>data_im_out(528),
            data_im_out(17)=>data_im_out(560),
            data_im_out(18)=>data_im_out(592),
            data_im_out(19)=>data_im_out(624),
            data_im_out(20)=>data_im_out(656),
            data_im_out(21)=>data_im_out(688),
            data_im_out(22)=>data_im_out(720),
            data_im_out(23)=>data_im_out(752),
            data_im_out(24)=>data_im_out(784),
            data_im_out(25)=>data_im_out(816),
            data_im_out(26)=>data_im_out(848),
            data_im_out(27)=>data_im_out(880),
            data_im_out(28)=>data_im_out(912),
            data_im_out(29)=>data_im_out(944),
            data_im_out(30)=>data_im_out(976),
            data_im_out(31)=>data_im_out(1008),
            data_im_out(32)=>data_im_out(1040),
            data_im_out(33)=>data_im_out(1072),
            data_im_out(34)=>data_im_out(1104),
            data_im_out(35)=>data_im_out(1136),
            data_im_out(36)=>data_im_out(1168),
            data_im_out(37)=>data_im_out(1200),
            data_im_out(38)=>data_im_out(1232),
            data_im_out(39)=>data_im_out(1264),
            data_im_out(40)=>data_im_out(1296),
            data_im_out(41)=>data_im_out(1328),
            data_im_out(42)=>data_im_out(1360),
            data_im_out(43)=>data_im_out(1392),
            data_im_out(44)=>data_im_out(1424),
            data_im_out(45)=>data_im_out(1456),
            data_im_out(46)=>data_im_out(1488),
            data_im_out(47)=>data_im_out(1520),
            data_im_out(48)=>data_im_out(1552),
            data_im_out(49)=>data_im_out(1584),
            data_im_out(50)=>data_im_out(1616),
            data_im_out(51)=>data_im_out(1648),
            data_im_out(52)=>data_im_out(1680),
            data_im_out(53)=>data_im_out(1712),
            data_im_out(54)=>data_im_out(1744),
            data_im_out(55)=>data_im_out(1776),
            data_im_out(56)=>data_im_out(1808),
            data_im_out(57)=>data_im_out(1840),
            data_im_out(58)=>data_im_out(1872),
            data_im_out(59)=>data_im_out(1904),
            data_im_out(60)=>data_im_out(1936),
            data_im_out(61)=>data_im_out(1968),
            data_im_out(62)=>data_im_out(2000),
            data_im_out(63)=>data_im_out(2032)
        );           

    URFFT_PT64_17 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(17),
            data_re_in(1)=>mul_re_out(49),
            data_re_in(2)=>mul_re_out(81),
            data_re_in(3)=>mul_re_out(113),
            data_re_in(4)=>mul_re_out(145),
            data_re_in(5)=>mul_re_out(177),
            data_re_in(6)=>mul_re_out(209),
            data_re_in(7)=>mul_re_out(241),
            data_re_in(8)=>mul_re_out(273),
            data_re_in(9)=>mul_re_out(305),
            data_re_in(10)=>mul_re_out(337),
            data_re_in(11)=>mul_re_out(369),
            data_re_in(12)=>mul_re_out(401),
            data_re_in(13)=>mul_re_out(433),
            data_re_in(14)=>mul_re_out(465),
            data_re_in(15)=>mul_re_out(497),
            data_re_in(16)=>mul_re_out(529),
            data_re_in(17)=>mul_re_out(561),
            data_re_in(18)=>mul_re_out(593),
            data_re_in(19)=>mul_re_out(625),
            data_re_in(20)=>mul_re_out(657),
            data_re_in(21)=>mul_re_out(689),
            data_re_in(22)=>mul_re_out(721),
            data_re_in(23)=>mul_re_out(753),
            data_re_in(24)=>mul_re_out(785),
            data_re_in(25)=>mul_re_out(817),
            data_re_in(26)=>mul_re_out(849),
            data_re_in(27)=>mul_re_out(881),
            data_re_in(28)=>mul_re_out(913),
            data_re_in(29)=>mul_re_out(945),
            data_re_in(30)=>mul_re_out(977),
            data_re_in(31)=>mul_re_out(1009),
            data_re_in(32)=>mul_re_out(1041),
            data_re_in(33)=>mul_re_out(1073),
            data_re_in(34)=>mul_re_out(1105),
            data_re_in(35)=>mul_re_out(1137),
            data_re_in(36)=>mul_re_out(1169),
            data_re_in(37)=>mul_re_out(1201),
            data_re_in(38)=>mul_re_out(1233),
            data_re_in(39)=>mul_re_out(1265),
            data_re_in(40)=>mul_re_out(1297),
            data_re_in(41)=>mul_re_out(1329),
            data_re_in(42)=>mul_re_out(1361),
            data_re_in(43)=>mul_re_out(1393),
            data_re_in(44)=>mul_re_out(1425),
            data_re_in(45)=>mul_re_out(1457),
            data_re_in(46)=>mul_re_out(1489),
            data_re_in(47)=>mul_re_out(1521),
            data_re_in(48)=>mul_re_out(1553),
            data_re_in(49)=>mul_re_out(1585),
            data_re_in(50)=>mul_re_out(1617),
            data_re_in(51)=>mul_re_out(1649),
            data_re_in(52)=>mul_re_out(1681),
            data_re_in(53)=>mul_re_out(1713),
            data_re_in(54)=>mul_re_out(1745),
            data_re_in(55)=>mul_re_out(1777),
            data_re_in(56)=>mul_re_out(1809),
            data_re_in(57)=>mul_re_out(1841),
            data_re_in(58)=>mul_re_out(1873),
            data_re_in(59)=>mul_re_out(1905),
            data_re_in(60)=>mul_re_out(1937),
            data_re_in(61)=>mul_re_out(1969),
            data_re_in(62)=>mul_re_out(2001),
            data_re_in(63)=>mul_re_out(2033),
            data_im_in(0)=>mul_im_out(17),
            data_im_in(1)=>mul_im_out(49),
            data_im_in(2)=>mul_im_out(81),
            data_im_in(3)=>mul_im_out(113),
            data_im_in(4)=>mul_im_out(145),
            data_im_in(5)=>mul_im_out(177),
            data_im_in(6)=>mul_im_out(209),
            data_im_in(7)=>mul_im_out(241),
            data_im_in(8)=>mul_im_out(273),
            data_im_in(9)=>mul_im_out(305),
            data_im_in(10)=>mul_im_out(337),
            data_im_in(11)=>mul_im_out(369),
            data_im_in(12)=>mul_im_out(401),
            data_im_in(13)=>mul_im_out(433),
            data_im_in(14)=>mul_im_out(465),
            data_im_in(15)=>mul_im_out(497),
            data_im_in(16)=>mul_im_out(529),
            data_im_in(17)=>mul_im_out(561),
            data_im_in(18)=>mul_im_out(593),
            data_im_in(19)=>mul_im_out(625),
            data_im_in(20)=>mul_im_out(657),
            data_im_in(21)=>mul_im_out(689),
            data_im_in(22)=>mul_im_out(721),
            data_im_in(23)=>mul_im_out(753),
            data_im_in(24)=>mul_im_out(785),
            data_im_in(25)=>mul_im_out(817),
            data_im_in(26)=>mul_im_out(849),
            data_im_in(27)=>mul_im_out(881),
            data_im_in(28)=>mul_im_out(913),
            data_im_in(29)=>mul_im_out(945),
            data_im_in(30)=>mul_im_out(977),
            data_im_in(31)=>mul_im_out(1009),
            data_im_in(32)=>mul_im_out(1041),
            data_im_in(33)=>mul_im_out(1073),
            data_im_in(34)=>mul_im_out(1105),
            data_im_in(35)=>mul_im_out(1137),
            data_im_in(36)=>mul_im_out(1169),
            data_im_in(37)=>mul_im_out(1201),
            data_im_in(38)=>mul_im_out(1233),
            data_im_in(39)=>mul_im_out(1265),
            data_im_in(40)=>mul_im_out(1297),
            data_im_in(41)=>mul_im_out(1329),
            data_im_in(42)=>mul_im_out(1361),
            data_im_in(43)=>mul_im_out(1393),
            data_im_in(44)=>mul_im_out(1425),
            data_im_in(45)=>mul_im_out(1457),
            data_im_in(46)=>mul_im_out(1489),
            data_im_in(47)=>mul_im_out(1521),
            data_im_in(48)=>mul_im_out(1553),
            data_im_in(49)=>mul_im_out(1585),
            data_im_in(50)=>mul_im_out(1617),
            data_im_in(51)=>mul_im_out(1649),
            data_im_in(52)=>mul_im_out(1681),
            data_im_in(53)=>mul_im_out(1713),
            data_im_in(54)=>mul_im_out(1745),
            data_im_in(55)=>mul_im_out(1777),
            data_im_in(56)=>mul_im_out(1809),
            data_im_in(57)=>mul_im_out(1841),
            data_im_in(58)=>mul_im_out(1873),
            data_im_in(59)=>mul_im_out(1905),
            data_im_in(60)=>mul_im_out(1937),
            data_im_in(61)=>mul_im_out(1969),
            data_im_in(62)=>mul_im_out(2001),
            data_im_in(63)=>mul_im_out(2033),
            data_re_out(0)=>data_re_out(17),
            data_re_out(1)=>data_re_out(49),
            data_re_out(2)=>data_re_out(81),
            data_re_out(3)=>data_re_out(113),
            data_re_out(4)=>data_re_out(145),
            data_re_out(5)=>data_re_out(177),
            data_re_out(6)=>data_re_out(209),
            data_re_out(7)=>data_re_out(241),
            data_re_out(8)=>data_re_out(273),
            data_re_out(9)=>data_re_out(305),
            data_re_out(10)=>data_re_out(337),
            data_re_out(11)=>data_re_out(369),
            data_re_out(12)=>data_re_out(401),
            data_re_out(13)=>data_re_out(433),
            data_re_out(14)=>data_re_out(465),
            data_re_out(15)=>data_re_out(497),
            data_re_out(16)=>data_re_out(529),
            data_re_out(17)=>data_re_out(561),
            data_re_out(18)=>data_re_out(593),
            data_re_out(19)=>data_re_out(625),
            data_re_out(20)=>data_re_out(657),
            data_re_out(21)=>data_re_out(689),
            data_re_out(22)=>data_re_out(721),
            data_re_out(23)=>data_re_out(753),
            data_re_out(24)=>data_re_out(785),
            data_re_out(25)=>data_re_out(817),
            data_re_out(26)=>data_re_out(849),
            data_re_out(27)=>data_re_out(881),
            data_re_out(28)=>data_re_out(913),
            data_re_out(29)=>data_re_out(945),
            data_re_out(30)=>data_re_out(977),
            data_re_out(31)=>data_re_out(1009),
            data_re_out(32)=>data_re_out(1041),
            data_re_out(33)=>data_re_out(1073),
            data_re_out(34)=>data_re_out(1105),
            data_re_out(35)=>data_re_out(1137),
            data_re_out(36)=>data_re_out(1169),
            data_re_out(37)=>data_re_out(1201),
            data_re_out(38)=>data_re_out(1233),
            data_re_out(39)=>data_re_out(1265),
            data_re_out(40)=>data_re_out(1297),
            data_re_out(41)=>data_re_out(1329),
            data_re_out(42)=>data_re_out(1361),
            data_re_out(43)=>data_re_out(1393),
            data_re_out(44)=>data_re_out(1425),
            data_re_out(45)=>data_re_out(1457),
            data_re_out(46)=>data_re_out(1489),
            data_re_out(47)=>data_re_out(1521),
            data_re_out(48)=>data_re_out(1553),
            data_re_out(49)=>data_re_out(1585),
            data_re_out(50)=>data_re_out(1617),
            data_re_out(51)=>data_re_out(1649),
            data_re_out(52)=>data_re_out(1681),
            data_re_out(53)=>data_re_out(1713),
            data_re_out(54)=>data_re_out(1745),
            data_re_out(55)=>data_re_out(1777),
            data_re_out(56)=>data_re_out(1809),
            data_re_out(57)=>data_re_out(1841),
            data_re_out(58)=>data_re_out(1873),
            data_re_out(59)=>data_re_out(1905),
            data_re_out(60)=>data_re_out(1937),
            data_re_out(61)=>data_re_out(1969),
            data_re_out(62)=>data_re_out(2001),
            data_re_out(63)=>data_re_out(2033),
            data_im_out(0)=>data_im_out(17),
            data_im_out(1)=>data_im_out(49),
            data_im_out(2)=>data_im_out(81),
            data_im_out(3)=>data_im_out(113),
            data_im_out(4)=>data_im_out(145),
            data_im_out(5)=>data_im_out(177),
            data_im_out(6)=>data_im_out(209),
            data_im_out(7)=>data_im_out(241),
            data_im_out(8)=>data_im_out(273),
            data_im_out(9)=>data_im_out(305),
            data_im_out(10)=>data_im_out(337),
            data_im_out(11)=>data_im_out(369),
            data_im_out(12)=>data_im_out(401),
            data_im_out(13)=>data_im_out(433),
            data_im_out(14)=>data_im_out(465),
            data_im_out(15)=>data_im_out(497),
            data_im_out(16)=>data_im_out(529),
            data_im_out(17)=>data_im_out(561),
            data_im_out(18)=>data_im_out(593),
            data_im_out(19)=>data_im_out(625),
            data_im_out(20)=>data_im_out(657),
            data_im_out(21)=>data_im_out(689),
            data_im_out(22)=>data_im_out(721),
            data_im_out(23)=>data_im_out(753),
            data_im_out(24)=>data_im_out(785),
            data_im_out(25)=>data_im_out(817),
            data_im_out(26)=>data_im_out(849),
            data_im_out(27)=>data_im_out(881),
            data_im_out(28)=>data_im_out(913),
            data_im_out(29)=>data_im_out(945),
            data_im_out(30)=>data_im_out(977),
            data_im_out(31)=>data_im_out(1009),
            data_im_out(32)=>data_im_out(1041),
            data_im_out(33)=>data_im_out(1073),
            data_im_out(34)=>data_im_out(1105),
            data_im_out(35)=>data_im_out(1137),
            data_im_out(36)=>data_im_out(1169),
            data_im_out(37)=>data_im_out(1201),
            data_im_out(38)=>data_im_out(1233),
            data_im_out(39)=>data_im_out(1265),
            data_im_out(40)=>data_im_out(1297),
            data_im_out(41)=>data_im_out(1329),
            data_im_out(42)=>data_im_out(1361),
            data_im_out(43)=>data_im_out(1393),
            data_im_out(44)=>data_im_out(1425),
            data_im_out(45)=>data_im_out(1457),
            data_im_out(46)=>data_im_out(1489),
            data_im_out(47)=>data_im_out(1521),
            data_im_out(48)=>data_im_out(1553),
            data_im_out(49)=>data_im_out(1585),
            data_im_out(50)=>data_im_out(1617),
            data_im_out(51)=>data_im_out(1649),
            data_im_out(52)=>data_im_out(1681),
            data_im_out(53)=>data_im_out(1713),
            data_im_out(54)=>data_im_out(1745),
            data_im_out(55)=>data_im_out(1777),
            data_im_out(56)=>data_im_out(1809),
            data_im_out(57)=>data_im_out(1841),
            data_im_out(58)=>data_im_out(1873),
            data_im_out(59)=>data_im_out(1905),
            data_im_out(60)=>data_im_out(1937),
            data_im_out(61)=>data_im_out(1969),
            data_im_out(62)=>data_im_out(2001),
            data_im_out(63)=>data_im_out(2033)
        );           

    URFFT_PT64_18 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(18),
            data_re_in(1)=>mul_re_out(50),
            data_re_in(2)=>mul_re_out(82),
            data_re_in(3)=>mul_re_out(114),
            data_re_in(4)=>mul_re_out(146),
            data_re_in(5)=>mul_re_out(178),
            data_re_in(6)=>mul_re_out(210),
            data_re_in(7)=>mul_re_out(242),
            data_re_in(8)=>mul_re_out(274),
            data_re_in(9)=>mul_re_out(306),
            data_re_in(10)=>mul_re_out(338),
            data_re_in(11)=>mul_re_out(370),
            data_re_in(12)=>mul_re_out(402),
            data_re_in(13)=>mul_re_out(434),
            data_re_in(14)=>mul_re_out(466),
            data_re_in(15)=>mul_re_out(498),
            data_re_in(16)=>mul_re_out(530),
            data_re_in(17)=>mul_re_out(562),
            data_re_in(18)=>mul_re_out(594),
            data_re_in(19)=>mul_re_out(626),
            data_re_in(20)=>mul_re_out(658),
            data_re_in(21)=>mul_re_out(690),
            data_re_in(22)=>mul_re_out(722),
            data_re_in(23)=>mul_re_out(754),
            data_re_in(24)=>mul_re_out(786),
            data_re_in(25)=>mul_re_out(818),
            data_re_in(26)=>mul_re_out(850),
            data_re_in(27)=>mul_re_out(882),
            data_re_in(28)=>mul_re_out(914),
            data_re_in(29)=>mul_re_out(946),
            data_re_in(30)=>mul_re_out(978),
            data_re_in(31)=>mul_re_out(1010),
            data_re_in(32)=>mul_re_out(1042),
            data_re_in(33)=>mul_re_out(1074),
            data_re_in(34)=>mul_re_out(1106),
            data_re_in(35)=>mul_re_out(1138),
            data_re_in(36)=>mul_re_out(1170),
            data_re_in(37)=>mul_re_out(1202),
            data_re_in(38)=>mul_re_out(1234),
            data_re_in(39)=>mul_re_out(1266),
            data_re_in(40)=>mul_re_out(1298),
            data_re_in(41)=>mul_re_out(1330),
            data_re_in(42)=>mul_re_out(1362),
            data_re_in(43)=>mul_re_out(1394),
            data_re_in(44)=>mul_re_out(1426),
            data_re_in(45)=>mul_re_out(1458),
            data_re_in(46)=>mul_re_out(1490),
            data_re_in(47)=>mul_re_out(1522),
            data_re_in(48)=>mul_re_out(1554),
            data_re_in(49)=>mul_re_out(1586),
            data_re_in(50)=>mul_re_out(1618),
            data_re_in(51)=>mul_re_out(1650),
            data_re_in(52)=>mul_re_out(1682),
            data_re_in(53)=>mul_re_out(1714),
            data_re_in(54)=>mul_re_out(1746),
            data_re_in(55)=>mul_re_out(1778),
            data_re_in(56)=>mul_re_out(1810),
            data_re_in(57)=>mul_re_out(1842),
            data_re_in(58)=>mul_re_out(1874),
            data_re_in(59)=>mul_re_out(1906),
            data_re_in(60)=>mul_re_out(1938),
            data_re_in(61)=>mul_re_out(1970),
            data_re_in(62)=>mul_re_out(2002),
            data_re_in(63)=>mul_re_out(2034),
            data_im_in(0)=>mul_im_out(18),
            data_im_in(1)=>mul_im_out(50),
            data_im_in(2)=>mul_im_out(82),
            data_im_in(3)=>mul_im_out(114),
            data_im_in(4)=>mul_im_out(146),
            data_im_in(5)=>mul_im_out(178),
            data_im_in(6)=>mul_im_out(210),
            data_im_in(7)=>mul_im_out(242),
            data_im_in(8)=>mul_im_out(274),
            data_im_in(9)=>mul_im_out(306),
            data_im_in(10)=>mul_im_out(338),
            data_im_in(11)=>mul_im_out(370),
            data_im_in(12)=>mul_im_out(402),
            data_im_in(13)=>mul_im_out(434),
            data_im_in(14)=>mul_im_out(466),
            data_im_in(15)=>mul_im_out(498),
            data_im_in(16)=>mul_im_out(530),
            data_im_in(17)=>mul_im_out(562),
            data_im_in(18)=>mul_im_out(594),
            data_im_in(19)=>mul_im_out(626),
            data_im_in(20)=>mul_im_out(658),
            data_im_in(21)=>mul_im_out(690),
            data_im_in(22)=>mul_im_out(722),
            data_im_in(23)=>mul_im_out(754),
            data_im_in(24)=>mul_im_out(786),
            data_im_in(25)=>mul_im_out(818),
            data_im_in(26)=>mul_im_out(850),
            data_im_in(27)=>mul_im_out(882),
            data_im_in(28)=>mul_im_out(914),
            data_im_in(29)=>mul_im_out(946),
            data_im_in(30)=>mul_im_out(978),
            data_im_in(31)=>mul_im_out(1010),
            data_im_in(32)=>mul_im_out(1042),
            data_im_in(33)=>mul_im_out(1074),
            data_im_in(34)=>mul_im_out(1106),
            data_im_in(35)=>mul_im_out(1138),
            data_im_in(36)=>mul_im_out(1170),
            data_im_in(37)=>mul_im_out(1202),
            data_im_in(38)=>mul_im_out(1234),
            data_im_in(39)=>mul_im_out(1266),
            data_im_in(40)=>mul_im_out(1298),
            data_im_in(41)=>mul_im_out(1330),
            data_im_in(42)=>mul_im_out(1362),
            data_im_in(43)=>mul_im_out(1394),
            data_im_in(44)=>mul_im_out(1426),
            data_im_in(45)=>mul_im_out(1458),
            data_im_in(46)=>mul_im_out(1490),
            data_im_in(47)=>mul_im_out(1522),
            data_im_in(48)=>mul_im_out(1554),
            data_im_in(49)=>mul_im_out(1586),
            data_im_in(50)=>mul_im_out(1618),
            data_im_in(51)=>mul_im_out(1650),
            data_im_in(52)=>mul_im_out(1682),
            data_im_in(53)=>mul_im_out(1714),
            data_im_in(54)=>mul_im_out(1746),
            data_im_in(55)=>mul_im_out(1778),
            data_im_in(56)=>mul_im_out(1810),
            data_im_in(57)=>mul_im_out(1842),
            data_im_in(58)=>mul_im_out(1874),
            data_im_in(59)=>mul_im_out(1906),
            data_im_in(60)=>mul_im_out(1938),
            data_im_in(61)=>mul_im_out(1970),
            data_im_in(62)=>mul_im_out(2002),
            data_im_in(63)=>mul_im_out(2034),
            data_re_out(0)=>data_re_out(18),
            data_re_out(1)=>data_re_out(50),
            data_re_out(2)=>data_re_out(82),
            data_re_out(3)=>data_re_out(114),
            data_re_out(4)=>data_re_out(146),
            data_re_out(5)=>data_re_out(178),
            data_re_out(6)=>data_re_out(210),
            data_re_out(7)=>data_re_out(242),
            data_re_out(8)=>data_re_out(274),
            data_re_out(9)=>data_re_out(306),
            data_re_out(10)=>data_re_out(338),
            data_re_out(11)=>data_re_out(370),
            data_re_out(12)=>data_re_out(402),
            data_re_out(13)=>data_re_out(434),
            data_re_out(14)=>data_re_out(466),
            data_re_out(15)=>data_re_out(498),
            data_re_out(16)=>data_re_out(530),
            data_re_out(17)=>data_re_out(562),
            data_re_out(18)=>data_re_out(594),
            data_re_out(19)=>data_re_out(626),
            data_re_out(20)=>data_re_out(658),
            data_re_out(21)=>data_re_out(690),
            data_re_out(22)=>data_re_out(722),
            data_re_out(23)=>data_re_out(754),
            data_re_out(24)=>data_re_out(786),
            data_re_out(25)=>data_re_out(818),
            data_re_out(26)=>data_re_out(850),
            data_re_out(27)=>data_re_out(882),
            data_re_out(28)=>data_re_out(914),
            data_re_out(29)=>data_re_out(946),
            data_re_out(30)=>data_re_out(978),
            data_re_out(31)=>data_re_out(1010),
            data_re_out(32)=>data_re_out(1042),
            data_re_out(33)=>data_re_out(1074),
            data_re_out(34)=>data_re_out(1106),
            data_re_out(35)=>data_re_out(1138),
            data_re_out(36)=>data_re_out(1170),
            data_re_out(37)=>data_re_out(1202),
            data_re_out(38)=>data_re_out(1234),
            data_re_out(39)=>data_re_out(1266),
            data_re_out(40)=>data_re_out(1298),
            data_re_out(41)=>data_re_out(1330),
            data_re_out(42)=>data_re_out(1362),
            data_re_out(43)=>data_re_out(1394),
            data_re_out(44)=>data_re_out(1426),
            data_re_out(45)=>data_re_out(1458),
            data_re_out(46)=>data_re_out(1490),
            data_re_out(47)=>data_re_out(1522),
            data_re_out(48)=>data_re_out(1554),
            data_re_out(49)=>data_re_out(1586),
            data_re_out(50)=>data_re_out(1618),
            data_re_out(51)=>data_re_out(1650),
            data_re_out(52)=>data_re_out(1682),
            data_re_out(53)=>data_re_out(1714),
            data_re_out(54)=>data_re_out(1746),
            data_re_out(55)=>data_re_out(1778),
            data_re_out(56)=>data_re_out(1810),
            data_re_out(57)=>data_re_out(1842),
            data_re_out(58)=>data_re_out(1874),
            data_re_out(59)=>data_re_out(1906),
            data_re_out(60)=>data_re_out(1938),
            data_re_out(61)=>data_re_out(1970),
            data_re_out(62)=>data_re_out(2002),
            data_re_out(63)=>data_re_out(2034),
            data_im_out(0)=>data_im_out(18),
            data_im_out(1)=>data_im_out(50),
            data_im_out(2)=>data_im_out(82),
            data_im_out(3)=>data_im_out(114),
            data_im_out(4)=>data_im_out(146),
            data_im_out(5)=>data_im_out(178),
            data_im_out(6)=>data_im_out(210),
            data_im_out(7)=>data_im_out(242),
            data_im_out(8)=>data_im_out(274),
            data_im_out(9)=>data_im_out(306),
            data_im_out(10)=>data_im_out(338),
            data_im_out(11)=>data_im_out(370),
            data_im_out(12)=>data_im_out(402),
            data_im_out(13)=>data_im_out(434),
            data_im_out(14)=>data_im_out(466),
            data_im_out(15)=>data_im_out(498),
            data_im_out(16)=>data_im_out(530),
            data_im_out(17)=>data_im_out(562),
            data_im_out(18)=>data_im_out(594),
            data_im_out(19)=>data_im_out(626),
            data_im_out(20)=>data_im_out(658),
            data_im_out(21)=>data_im_out(690),
            data_im_out(22)=>data_im_out(722),
            data_im_out(23)=>data_im_out(754),
            data_im_out(24)=>data_im_out(786),
            data_im_out(25)=>data_im_out(818),
            data_im_out(26)=>data_im_out(850),
            data_im_out(27)=>data_im_out(882),
            data_im_out(28)=>data_im_out(914),
            data_im_out(29)=>data_im_out(946),
            data_im_out(30)=>data_im_out(978),
            data_im_out(31)=>data_im_out(1010),
            data_im_out(32)=>data_im_out(1042),
            data_im_out(33)=>data_im_out(1074),
            data_im_out(34)=>data_im_out(1106),
            data_im_out(35)=>data_im_out(1138),
            data_im_out(36)=>data_im_out(1170),
            data_im_out(37)=>data_im_out(1202),
            data_im_out(38)=>data_im_out(1234),
            data_im_out(39)=>data_im_out(1266),
            data_im_out(40)=>data_im_out(1298),
            data_im_out(41)=>data_im_out(1330),
            data_im_out(42)=>data_im_out(1362),
            data_im_out(43)=>data_im_out(1394),
            data_im_out(44)=>data_im_out(1426),
            data_im_out(45)=>data_im_out(1458),
            data_im_out(46)=>data_im_out(1490),
            data_im_out(47)=>data_im_out(1522),
            data_im_out(48)=>data_im_out(1554),
            data_im_out(49)=>data_im_out(1586),
            data_im_out(50)=>data_im_out(1618),
            data_im_out(51)=>data_im_out(1650),
            data_im_out(52)=>data_im_out(1682),
            data_im_out(53)=>data_im_out(1714),
            data_im_out(54)=>data_im_out(1746),
            data_im_out(55)=>data_im_out(1778),
            data_im_out(56)=>data_im_out(1810),
            data_im_out(57)=>data_im_out(1842),
            data_im_out(58)=>data_im_out(1874),
            data_im_out(59)=>data_im_out(1906),
            data_im_out(60)=>data_im_out(1938),
            data_im_out(61)=>data_im_out(1970),
            data_im_out(62)=>data_im_out(2002),
            data_im_out(63)=>data_im_out(2034)
        );           

    URFFT_PT64_19 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(19),
            data_re_in(1)=>mul_re_out(51),
            data_re_in(2)=>mul_re_out(83),
            data_re_in(3)=>mul_re_out(115),
            data_re_in(4)=>mul_re_out(147),
            data_re_in(5)=>mul_re_out(179),
            data_re_in(6)=>mul_re_out(211),
            data_re_in(7)=>mul_re_out(243),
            data_re_in(8)=>mul_re_out(275),
            data_re_in(9)=>mul_re_out(307),
            data_re_in(10)=>mul_re_out(339),
            data_re_in(11)=>mul_re_out(371),
            data_re_in(12)=>mul_re_out(403),
            data_re_in(13)=>mul_re_out(435),
            data_re_in(14)=>mul_re_out(467),
            data_re_in(15)=>mul_re_out(499),
            data_re_in(16)=>mul_re_out(531),
            data_re_in(17)=>mul_re_out(563),
            data_re_in(18)=>mul_re_out(595),
            data_re_in(19)=>mul_re_out(627),
            data_re_in(20)=>mul_re_out(659),
            data_re_in(21)=>mul_re_out(691),
            data_re_in(22)=>mul_re_out(723),
            data_re_in(23)=>mul_re_out(755),
            data_re_in(24)=>mul_re_out(787),
            data_re_in(25)=>mul_re_out(819),
            data_re_in(26)=>mul_re_out(851),
            data_re_in(27)=>mul_re_out(883),
            data_re_in(28)=>mul_re_out(915),
            data_re_in(29)=>mul_re_out(947),
            data_re_in(30)=>mul_re_out(979),
            data_re_in(31)=>mul_re_out(1011),
            data_re_in(32)=>mul_re_out(1043),
            data_re_in(33)=>mul_re_out(1075),
            data_re_in(34)=>mul_re_out(1107),
            data_re_in(35)=>mul_re_out(1139),
            data_re_in(36)=>mul_re_out(1171),
            data_re_in(37)=>mul_re_out(1203),
            data_re_in(38)=>mul_re_out(1235),
            data_re_in(39)=>mul_re_out(1267),
            data_re_in(40)=>mul_re_out(1299),
            data_re_in(41)=>mul_re_out(1331),
            data_re_in(42)=>mul_re_out(1363),
            data_re_in(43)=>mul_re_out(1395),
            data_re_in(44)=>mul_re_out(1427),
            data_re_in(45)=>mul_re_out(1459),
            data_re_in(46)=>mul_re_out(1491),
            data_re_in(47)=>mul_re_out(1523),
            data_re_in(48)=>mul_re_out(1555),
            data_re_in(49)=>mul_re_out(1587),
            data_re_in(50)=>mul_re_out(1619),
            data_re_in(51)=>mul_re_out(1651),
            data_re_in(52)=>mul_re_out(1683),
            data_re_in(53)=>mul_re_out(1715),
            data_re_in(54)=>mul_re_out(1747),
            data_re_in(55)=>mul_re_out(1779),
            data_re_in(56)=>mul_re_out(1811),
            data_re_in(57)=>mul_re_out(1843),
            data_re_in(58)=>mul_re_out(1875),
            data_re_in(59)=>mul_re_out(1907),
            data_re_in(60)=>mul_re_out(1939),
            data_re_in(61)=>mul_re_out(1971),
            data_re_in(62)=>mul_re_out(2003),
            data_re_in(63)=>mul_re_out(2035),
            data_im_in(0)=>mul_im_out(19),
            data_im_in(1)=>mul_im_out(51),
            data_im_in(2)=>mul_im_out(83),
            data_im_in(3)=>mul_im_out(115),
            data_im_in(4)=>mul_im_out(147),
            data_im_in(5)=>mul_im_out(179),
            data_im_in(6)=>mul_im_out(211),
            data_im_in(7)=>mul_im_out(243),
            data_im_in(8)=>mul_im_out(275),
            data_im_in(9)=>mul_im_out(307),
            data_im_in(10)=>mul_im_out(339),
            data_im_in(11)=>mul_im_out(371),
            data_im_in(12)=>mul_im_out(403),
            data_im_in(13)=>mul_im_out(435),
            data_im_in(14)=>mul_im_out(467),
            data_im_in(15)=>mul_im_out(499),
            data_im_in(16)=>mul_im_out(531),
            data_im_in(17)=>mul_im_out(563),
            data_im_in(18)=>mul_im_out(595),
            data_im_in(19)=>mul_im_out(627),
            data_im_in(20)=>mul_im_out(659),
            data_im_in(21)=>mul_im_out(691),
            data_im_in(22)=>mul_im_out(723),
            data_im_in(23)=>mul_im_out(755),
            data_im_in(24)=>mul_im_out(787),
            data_im_in(25)=>mul_im_out(819),
            data_im_in(26)=>mul_im_out(851),
            data_im_in(27)=>mul_im_out(883),
            data_im_in(28)=>mul_im_out(915),
            data_im_in(29)=>mul_im_out(947),
            data_im_in(30)=>mul_im_out(979),
            data_im_in(31)=>mul_im_out(1011),
            data_im_in(32)=>mul_im_out(1043),
            data_im_in(33)=>mul_im_out(1075),
            data_im_in(34)=>mul_im_out(1107),
            data_im_in(35)=>mul_im_out(1139),
            data_im_in(36)=>mul_im_out(1171),
            data_im_in(37)=>mul_im_out(1203),
            data_im_in(38)=>mul_im_out(1235),
            data_im_in(39)=>mul_im_out(1267),
            data_im_in(40)=>mul_im_out(1299),
            data_im_in(41)=>mul_im_out(1331),
            data_im_in(42)=>mul_im_out(1363),
            data_im_in(43)=>mul_im_out(1395),
            data_im_in(44)=>mul_im_out(1427),
            data_im_in(45)=>mul_im_out(1459),
            data_im_in(46)=>mul_im_out(1491),
            data_im_in(47)=>mul_im_out(1523),
            data_im_in(48)=>mul_im_out(1555),
            data_im_in(49)=>mul_im_out(1587),
            data_im_in(50)=>mul_im_out(1619),
            data_im_in(51)=>mul_im_out(1651),
            data_im_in(52)=>mul_im_out(1683),
            data_im_in(53)=>mul_im_out(1715),
            data_im_in(54)=>mul_im_out(1747),
            data_im_in(55)=>mul_im_out(1779),
            data_im_in(56)=>mul_im_out(1811),
            data_im_in(57)=>mul_im_out(1843),
            data_im_in(58)=>mul_im_out(1875),
            data_im_in(59)=>mul_im_out(1907),
            data_im_in(60)=>mul_im_out(1939),
            data_im_in(61)=>mul_im_out(1971),
            data_im_in(62)=>mul_im_out(2003),
            data_im_in(63)=>mul_im_out(2035),
            data_re_out(0)=>data_re_out(19),
            data_re_out(1)=>data_re_out(51),
            data_re_out(2)=>data_re_out(83),
            data_re_out(3)=>data_re_out(115),
            data_re_out(4)=>data_re_out(147),
            data_re_out(5)=>data_re_out(179),
            data_re_out(6)=>data_re_out(211),
            data_re_out(7)=>data_re_out(243),
            data_re_out(8)=>data_re_out(275),
            data_re_out(9)=>data_re_out(307),
            data_re_out(10)=>data_re_out(339),
            data_re_out(11)=>data_re_out(371),
            data_re_out(12)=>data_re_out(403),
            data_re_out(13)=>data_re_out(435),
            data_re_out(14)=>data_re_out(467),
            data_re_out(15)=>data_re_out(499),
            data_re_out(16)=>data_re_out(531),
            data_re_out(17)=>data_re_out(563),
            data_re_out(18)=>data_re_out(595),
            data_re_out(19)=>data_re_out(627),
            data_re_out(20)=>data_re_out(659),
            data_re_out(21)=>data_re_out(691),
            data_re_out(22)=>data_re_out(723),
            data_re_out(23)=>data_re_out(755),
            data_re_out(24)=>data_re_out(787),
            data_re_out(25)=>data_re_out(819),
            data_re_out(26)=>data_re_out(851),
            data_re_out(27)=>data_re_out(883),
            data_re_out(28)=>data_re_out(915),
            data_re_out(29)=>data_re_out(947),
            data_re_out(30)=>data_re_out(979),
            data_re_out(31)=>data_re_out(1011),
            data_re_out(32)=>data_re_out(1043),
            data_re_out(33)=>data_re_out(1075),
            data_re_out(34)=>data_re_out(1107),
            data_re_out(35)=>data_re_out(1139),
            data_re_out(36)=>data_re_out(1171),
            data_re_out(37)=>data_re_out(1203),
            data_re_out(38)=>data_re_out(1235),
            data_re_out(39)=>data_re_out(1267),
            data_re_out(40)=>data_re_out(1299),
            data_re_out(41)=>data_re_out(1331),
            data_re_out(42)=>data_re_out(1363),
            data_re_out(43)=>data_re_out(1395),
            data_re_out(44)=>data_re_out(1427),
            data_re_out(45)=>data_re_out(1459),
            data_re_out(46)=>data_re_out(1491),
            data_re_out(47)=>data_re_out(1523),
            data_re_out(48)=>data_re_out(1555),
            data_re_out(49)=>data_re_out(1587),
            data_re_out(50)=>data_re_out(1619),
            data_re_out(51)=>data_re_out(1651),
            data_re_out(52)=>data_re_out(1683),
            data_re_out(53)=>data_re_out(1715),
            data_re_out(54)=>data_re_out(1747),
            data_re_out(55)=>data_re_out(1779),
            data_re_out(56)=>data_re_out(1811),
            data_re_out(57)=>data_re_out(1843),
            data_re_out(58)=>data_re_out(1875),
            data_re_out(59)=>data_re_out(1907),
            data_re_out(60)=>data_re_out(1939),
            data_re_out(61)=>data_re_out(1971),
            data_re_out(62)=>data_re_out(2003),
            data_re_out(63)=>data_re_out(2035),
            data_im_out(0)=>data_im_out(19),
            data_im_out(1)=>data_im_out(51),
            data_im_out(2)=>data_im_out(83),
            data_im_out(3)=>data_im_out(115),
            data_im_out(4)=>data_im_out(147),
            data_im_out(5)=>data_im_out(179),
            data_im_out(6)=>data_im_out(211),
            data_im_out(7)=>data_im_out(243),
            data_im_out(8)=>data_im_out(275),
            data_im_out(9)=>data_im_out(307),
            data_im_out(10)=>data_im_out(339),
            data_im_out(11)=>data_im_out(371),
            data_im_out(12)=>data_im_out(403),
            data_im_out(13)=>data_im_out(435),
            data_im_out(14)=>data_im_out(467),
            data_im_out(15)=>data_im_out(499),
            data_im_out(16)=>data_im_out(531),
            data_im_out(17)=>data_im_out(563),
            data_im_out(18)=>data_im_out(595),
            data_im_out(19)=>data_im_out(627),
            data_im_out(20)=>data_im_out(659),
            data_im_out(21)=>data_im_out(691),
            data_im_out(22)=>data_im_out(723),
            data_im_out(23)=>data_im_out(755),
            data_im_out(24)=>data_im_out(787),
            data_im_out(25)=>data_im_out(819),
            data_im_out(26)=>data_im_out(851),
            data_im_out(27)=>data_im_out(883),
            data_im_out(28)=>data_im_out(915),
            data_im_out(29)=>data_im_out(947),
            data_im_out(30)=>data_im_out(979),
            data_im_out(31)=>data_im_out(1011),
            data_im_out(32)=>data_im_out(1043),
            data_im_out(33)=>data_im_out(1075),
            data_im_out(34)=>data_im_out(1107),
            data_im_out(35)=>data_im_out(1139),
            data_im_out(36)=>data_im_out(1171),
            data_im_out(37)=>data_im_out(1203),
            data_im_out(38)=>data_im_out(1235),
            data_im_out(39)=>data_im_out(1267),
            data_im_out(40)=>data_im_out(1299),
            data_im_out(41)=>data_im_out(1331),
            data_im_out(42)=>data_im_out(1363),
            data_im_out(43)=>data_im_out(1395),
            data_im_out(44)=>data_im_out(1427),
            data_im_out(45)=>data_im_out(1459),
            data_im_out(46)=>data_im_out(1491),
            data_im_out(47)=>data_im_out(1523),
            data_im_out(48)=>data_im_out(1555),
            data_im_out(49)=>data_im_out(1587),
            data_im_out(50)=>data_im_out(1619),
            data_im_out(51)=>data_im_out(1651),
            data_im_out(52)=>data_im_out(1683),
            data_im_out(53)=>data_im_out(1715),
            data_im_out(54)=>data_im_out(1747),
            data_im_out(55)=>data_im_out(1779),
            data_im_out(56)=>data_im_out(1811),
            data_im_out(57)=>data_im_out(1843),
            data_im_out(58)=>data_im_out(1875),
            data_im_out(59)=>data_im_out(1907),
            data_im_out(60)=>data_im_out(1939),
            data_im_out(61)=>data_im_out(1971),
            data_im_out(62)=>data_im_out(2003),
            data_im_out(63)=>data_im_out(2035)
        );           

    URFFT_PT64_20 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(20),
            data_re_in(1)=>mul_re_out(52),
            data_re_in(2)=>mul_re_out(84),
            data_re_in(3)=>mul_re_out(116),
            data_re_in(4)=>mul_re_out(148),
            data_re_in(5)=>mul_re_out(180),
            data_re_in(6)=>mul_re_out(212),
            data_re_in(7)=>mul_re_out(244),
            data_re_in(8)=>mul_re_out(276),
            data_re_in(9)=>mul_re_out(308),
            data_re_in(10)=>mul_re_out(340),
            data_re_in(11)=>mul_re_out(372),
            data_re_in(12)=>mul_re_out(404),
            data_re_in(13)=>mul_re_out(436),
            data_re_in(14)=>mul_re_out(468),
            data_re_in(15)=>mul_re_out(500),
            data_re_in(16)=>mul_re_out(532),
            data_re_in(17)=>mul_re_out(564),
            data_re_in(18)=>mul_re_out(596),
            data_re_in(19)=>mul_re_out(628),
            data_re_in(20)=>mul_re_out(660),
            data_re_in(21)=>mul_re_out(692),
            data_re_in(22)=>mul_re_out(724),
            data_re_in(23)=>mul_re_out(756),
            data_re_in(24)=>mul_re_out(788),
            data_re_in(25)=>mul_re_out(820),
            data_re_in(26)=>mul_re_out(852),
            data_re_in(27)=>mul_re_out(884),
            data_re_in(28)=>mul_re_out(916),
            data_re_in(29)=>mul_re_out(948),
            data_re_in(30)=>mul_re_out(980),
            data_re_in(31)=>mul_re_out(1012),
            data_re_in(32)=>mul_re_out(1044),
            data_re_in(33)=>mul_re_out(1076),
            data_re_in(34)=>mul_re_out(1108),
            data_re_in(35)=>mul_re_out(1140),
            data_re_in(36)=>mul_re_out(1172),
            data_re_in(37)=>mul_re_out(1204),
            data_re_in(38)=>mul_re_out(1236),
            data_re_in(39)=>mul_re_out(1268),
            data_re_in(40)=>mul_re_out(1300),
            data_re_in(41)=>mul_re_out(1332),
            data_re_in(42)=>mul_re_out(1364),
            data_re_in(43)=>mul_re_out(1396),
            data_re_in(44)=>mul_re_out(1428),
            data_re_in(45)=>mul_re_out(1460),
            data_re_in(46)=>mul_re_out(1492),
            data_re_in(47)=>mul_re_out(1524),
            data_re_in(48)=>mul_re_out(1556),
            data_re_in(49)=>mul_re_out(1588),
            data_re_in(50)=>mul_re_out(1620),
            data_re_in(51)=>mul_re_out(1652),
            data_re_in(52)=>mul_re_out(1684),
            data_re_in(53)=>mul_re_out(1716),
            data_re_in(54)=>mul_re_out(1748),
            data_re_in(55)=>mul_re_out(1780),
            data_re_in(56)=>mul_re_out(1812),
            data_re_in(57)=>mul_re_out(1844),
            data_re_in(58)=>mul_re_out(1876),
            data_re_in(59)=>mul_re_out(1908),
            data_re_in(60)=>mul_re_out(1940),
            data_re_in(61)=>mul_re_out(1972),
            data_re_in(62)=>mul_re_out(2004),
            data_re_in(63)=>mul_re_out(2036),
            data_im_in(0)=>mul_im_out(20),
            data_im_in(1)=>mul_im_out(52),
            data_im_in(2)=>mul_im_out(84),
            data_im_in(3)=>mul_im_out(116),
            data_im_in(4)=>mul_im_out(148),
            data_im_in(5)=>mul_im_out(180),
            data_im_in(6)=>mul_im_out(212),
            data_im_in(7)=>mul_im_out(244),
            data_im_in(8)=>mul_im_out(276),
            data_im_in(9)=>mul_im_out(308),
            data_im_in(10)=>mul_im_out(340),
            data_im_in(11)=>mul_im_out(372),
            data_im_in(12)=>mul_im_out(404),
            data_im_in(13)=>mul_im_out(436),
            data_im_in(14)=>mul_im_out(468),
            data_im_in(15)=>mul_im_out(500),
            data_im_in(16)=>mul_im_out(532),
            data_im_in(17)=>mul_im_out(564),
            data_im_in(18)=>mul_im_out(596),
            data_im_in(19)=>mul_im_out(628),
            data_im_in(20)=>mul_im_out(660),
            data_im_in(21)=>mul_im_out(692),
            data_im_in(22)=>mul_im_out(724),
            data_im_in(23)=>mul_im_out(756),
            data_im_in(24)=>mul_im_out(788),
            data_im_in(25)=>mul_im_out(820),
            data_im_in(26)=>mul_im_out(852),
            data_im_in(27)=>mul_im_out(884),
            data_im_in(28)=>mul_im_out(916),
            data_im_in(29)=>mul_im_out(948),
            data_im_in(30)=>mul_im_out(980),
            data_im_in(31)=>mul_im_out(1012),
            data_im_in(32)=>mul_im_out(1044),
            data_im_in(33)=>mul_im_out(1076),
            data_im_in(34)=>mul_im_out(1108),
            data_im_in(35)=>mul_im_out(1140),
            data_im_in(36)=>mul_im_out(1172),
            data_im_in(37)=>mul_im_out(1204),
            data_im_in(38)=>mul_im_out(1236),
            data_im_in(39)=>mul_im_out(1268),
            data_im_in(40)=>mul_im_out(1300),
            data_im_in(41)=>mul_im_out(1332),
            data_im_in(42)=>mul_im_out(1364),
            data_im_in(43)=>mul_im_out(1396),
            data_im_in(44)=>mul_im_out(1428),
            data_im_in(45)=>mul_im_out(1460),
            data_im_in(46)=>mul_im_out(1492),
            data_im_in(47)=>mul_im_out(1524),
            data_im_in(48)=>mul_im_out(1556),
            data_im_in(49)=>mul_im_out(1588),
            data_im_in(50)=>mul_im_out(1620),
            data_im_in(51)=>mul_im_out(1652),
            data_im_in(52)=>mul_im_out(1684),
            data_im_in(53)=>mul_im_out(1716),
            data_im_in(54)=>mul_im_out(1748),
            data_im_in(55)=>mul_im_out(1780),
            data_im_in(56)=>mul_im_out(1812),
            data_im_in(57)=>mul_im_out(1844),
            data_im_in(58)=>mul_im_out(1876),
            data_im_in(59)=>mul_im_out(1908),
            data_im_in(60)=>mul_im_out(1940),
            data_im_in(61)=>mul_im_out(1972),
            data_im_in(62)=>mul_im_out(2004),
            data_im_in(63)=>mul_im_out(2036),
            data_re_out(0)=>data_re_out(20),
            data_re_out(1)=>data_re_out(52),
            data_re_out(2)=>data_re_out(84),
            data_re_out(3)=>data_re_out(116),
            data_re_out(4)=>data_re_out(148),
            data_re_out(5)=>data_re_out(180),
            data_re_out(6)=>data_re_out(212),
            data_re_out(7)=>data_re_out(244),
            data_re_out(8)=>data_re_out(276),
            data_re_out(9)=>data_re_out(308),
            data_re_out(10)=>data_re_out(340),
            data_re_out(11)=>data_re_out(372),
            data_re_out(12)=>data_re_out(404),
            data_re_out(13)=>data_re_out(436),
            data_re_out(14)=>data_re_out(468),
            data_re_out(15)=>data_re_out(500),
            data_re_out(16)=>data_re_out(532),
            data_re_out(17)=>data_re_out(564),
            data_re_out(18)=>data_re_out(596),
            data_re_out(19)=>data_re_out(628),
            data_re_out(20)=>data_re_out(660),
            data_re_out(21)=>data_re_out(692),
            data_re_out(22)=>data_re_out(724),
            data_re_out(23)=>data_re_out(756),
            data_re_out(24)=>data_re_out(788),
            data_re_out(25)=>data_re_out(820),
            data_re_out(26)=>data_re_out(852),
            data_re_out(27)=>data_re_out(884),
            data_re_out(28)=>data_re_out(916),
            data_re_out(29)=>data_re_out(948),
            data_re_out(30)=>data_re_out(980),
            data_re_out(31)=>data_re_out(1012),
            data_re_out(32)=>data_re_out(1044),
            data_re_out(33)=>data_re_out(1076),
            data_re_out(34)=>data_re_out(1108),
            data_re_out(35)=>data_re_out(1140),
            data_re_out(36)=>data_re_out(1172),
            data_re_out(37)=>data_re_out(1204),
            data_re_out(38)=>data_re_out(1236),
            data_re_out(39)=>data_re_out(1268),
            data_re_out(40)=>data_re_out(1300),
            data_re_out(41)=>data_re_out(1332),
            data_re_out(42)=>data_re_out(1364),
            data_re_out(43)=>data_re_out(1396),
            data_re_out(44)=>data_re_out(1428),
            data_re_out(45)=>data_re_out(1460),
            data_re_out(46)=>data_re_out(1492),
            data_re_out(47)=>data_re_out(1524),
            data_re_out(48)=>data_re_out(1556),
            data_re_out(49)=>data_re_out(1588),
            data_re_out(50)=>data_re_out(1620),
            data_re_out(51)=>data_re_out(1652),
            data_re_out(52)=>data_re_out(1684),
            data_re_out(53)=>data_re_out(1716),
            data_re_out(54)=>data_re_out(1748),
            data_re_out(55)=>data_re_out(1780),
            data_re_out(56)=>data_re_out(1812),
            data_re_out(57)=>data_re_out(1844),
            data_re_out(58)=>data_re_out(1876),
            data_re_out(59)=>data_re_out(1908),
            data_re_out(60)=>data_re_out(1940),
            data_re_out(61)=>data_re_out(1972),
            data_re_out(62)=>data_re_out(2004),
            data_re_out(63)=>data_re_out(2036),
            data_im_out(0)=>data_im_out(20),
            data_im_out(1)=>data_im_out(52),
            data_im_out(2)=>data_im_out(84),
            data_im_out(3)=>data_im_out(116),
            data_im_out(4)=>data_im_out(148),
            data_im_out(5)=>data_im_out(180),
            data_im_out(6)=>data_im_out(212),
            data_im_out(7)=>data_im_out(244),
            data_im_out(8)=>data_im_out(276),
            data_im_out(9)=>data_im_out(308),
            data_im_out(10)=>data_im_out(340),
            data_im_out(11)=>data_im_out(372),
            data_im_out(12)=>data_im_out(404),
            data_im_out(13)=>data_im_out(436),
            data_im_out(14)=>data_im_out(468),
            data_im_out(15)=>data_im_out(500),
            data_im_out(16)=>data_im_out(532),
            data_im_out(17)=>data_im_out(564),
            data_im_out(18)=>data_im_out(596),
            data_im_out(19)=>data_im_out(628),
            data_im_out(20)=>data_im_out(660),
            data_im_out(21)=>data_im_out(692),
            data_im_out(22)=>data_im_out(724),
            data_im_out(23)=>data_im_out(756),
            data_im_out(24)=>data_im_out(788),
            data_im_out(25)=>data_im_out(820),
            data_im_out(26)=>data_im_out(852),
            data_im_out(27)=>data_im_out(884),
            data_im_out(28)=>data_im_out(916),
            data_im_out(29)=>data_im_out(948),
            data_im_out(30)=>data_im_out(980),
            data_im_out(31)=>data_im_out(1012),
            data_im_out(32)=>data_im_out(1044),
            data_im_out(33)=>data_im_out(1076),
            data_im_out(34)=>data_im_out(1108),
            data_im_out(35)=>data_im_out(1140),
            data_im_out(36)=>data_im_out(1172),
            data_im_out(37)=>data_im_out(1204),
            data_im_out(38)=>data_im_out(1236),
            data_im_out(39)=>data_im_out(1268),
            data_im_out(40)=>data_im_out(1300),
            data_im_out(41)=>data_im_out(1332),
            data_im_out(42)=>data_im_out(1364),
            data_im_out(43)=>data_im_out(1396),
            data_im_out(44)=>data_im_out(1428),
            data_im_out(45)=>data_im_out(1460),
            data_im_out(46)=>data_im_out(1492),
            data_im_out(47)=>data_im_out(1524),
            data_im_out(48)=>data_im_out(1556),
            data_im_out(49)=>data_im_out(1588),
            data_im_out(50)=>data_im_out(1620),
            data_im_out(51)=>data_im_out(1652),
            data_im_out(52)=>data_im_out(1684),
            data_im_out(53)=>data_im_out(1716),
            data_im_out(54)=>data_im_out(1748),
            data_im_out(55)=>data_im_out(1780),
            data_im_out(56)=>data_im_out(1812),
            data_im_out(57)=>data_im_out(1844),
            data_im_out(58)=>data_im_out(1876),
            data_im_out(59)=>data_im_out(1908),
            data_im_out(60)=>data_im_out(1940),
            data_im_out(61)=>data_im_out(1972),
            data_im_out(62)=>data_im_out(2004),
            data_im_out(63)=>data_im_out(2036)
        );           

    URFFT_PT64_21 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(21),
            data_re_in(1)=>mul_re_out(53),
            data_re_in(2)=>mul_re_out(85),
            data_re_in(3)=>mul_re_out(117),
            data_re_in(4)=>mul_re_out(149),
            data_re_in(5)=>mul_re_out(181),
            data_re_in(6)=>mul_re_out(213),
            data_re_in(7)=>mul_re_out(245),
            data_re_in(8)=>mul_re_out(277),
            data_re_in(9)=>mul_re_out(309),
            data_re_in(10)=>mul_re_out(341),
            data_re_in(11)=>mul_re_out(373),
            data_re_in(12)=>mul_re_out(405),
            data_re_in(13)=>mul_re_out(437),
            data_re_in(14)=>mul_re_out(469),
            data_re_in(15)=>mul_re_out(501),
            data_re_in(16)=>mul_re_out(533),
            data_re_in(17)=>mul_re_out(565),
            data_re_in(18)=>mul_re_out(597),
            data_re_in(19)=>mul_re_out(629),
            data_re_in(20)=>mul_re_out(661),
            data_re_in(21)=>mul_re_out(693),
            data_re_in(22)=>mul_re_out(725),
            data_re_in(23)=>mul_re_out(757),
            data_re_in(24)=>mul_re_out(789),
            data_re_in(25)=>mul_re_out(821),
            data_re_in(26)=>mul_re_out(853),
            data_re_in(27)=>mul_re_out(885),
            data_re_in(28)=>mul_re_out(917),
            data_re_in(29)=>mul_re_out(949),
            data_re_in(30)=>mul_re_out(981),
            data_re_in(31)=>mul_re_out(1013),
            data_re_in(32)=>mul_re_out(1045),
            data_re_in(33)=>mul_re_out(1077),
            data_re_in(34)=>mul_re_out(1109),
            data_re_in(35)=>mul_re_out(1141),
            data_re_in(36)=>mul_re_out(1173),
            data_re_in(37)=>mul_re_out(1205),
            data_re_in(38)=>mul_re_out(1237),
            data_re_in(39)=>mul_re_out(1269),
            data_re_in(40)=>mul_re_out(1301),
            data_re_in(41)=>mul_re_out(1333),
            data_re_in(42)=>mul_re_out(1365),
            data_re_in(43)=>mul_re_out(1397),
            data_re_in(44)=>mul_re_out(1429),
            data_re_in(45)=>mul_re_out(1461),
            data_re_in(46)=>mul_re_out(1493),
            data_re_in(47)=>mul_re_out(1525),
            data_re_in(48)=>mul_re_out(1557),
            data_re_in(49)=>mul_re_out(1589),
            data_re_in(50)=>mul_re_out(1621),
            data_re_in(51)=>mul_re_out(1653),
            data_re_in(52)=>mul_re_out(1685),
            data_re_in(53)=>mul_re_out(1717),
            data_re_in(54)=>mul_re_out(1749),
            data_re_in(55)=>mul_re_out(1781),
            data_re_in(56)=>mul_re_out(1813),
            data_re_in(57)=>mul_re_out(1845),
            data_re_in(58)=>mul_re_out(1877),
            data_re_in(59)=>mul_re_out(1909),
            data_re_in(60)=>mul_re_out(1941),
            data_re_in(61)=>mul_re_out(1973),
            data_re_in(62)=>mul_re_out(2005),
            data_re_in(63)=>mul_re_out(2037),
            data_im_in(0)=>mul_im_out(21),
            data_im_in(1)=>mul_im_out(53),
            data_im_in(2)=>mul_im_out(85),
            data_im_in(3)=>mul_im_out(117),
            data_im_in(4)=>mul_im_out(149),
            data_im_in(5)=>mul_im_out(181),
            data_im_in(6)=>mul_im_out(213),
            data_im_in(7)=>mul_im_out(245),
            data_im_in(8)=>mul_im_out(277),
            data_im_in(9)=>mul_im_out(309),
            data_im_in(10)=>mul_im_out(341),
            data_im_in(11)=>mul_im_out(373),
            data_im_in(12)=>mul_im_out(405),
            data_im_in(13)=>mul_im_out(437),
            data_im_in(14)=>mul_im_out(469),
            data_im_in(15)=>mul_im_out(501),
            data_im_in(16)=>mul_im_out(533),
            data_im_in(17)=>mul_im_out(565),
            data_im_in(18)=>mul_im_out(597),
            data_im_in(19)=>mul_im_out(629),
            data_im_in(20)=>mul_im_out(661),
            data_im_in(21)=>mul_im_out(693),
            data_im_in(22)=>mul_im_out(725),
            data_im_in(23)=>mul_im_out(757),
            data_im_in(24)=>mul_im_out(789),
            data_im_in(25)=>mul_im_out(821),
            data_im_in(26)=>mul_im_out(853),
            data_im_in(27)=>mul_im_out(885),
            data_im_in(28)=>mul_im_out(917),
            data_im_in(29)=>mul_im_out(949),
            data_im_in(30)=>mul_im_out(981),
            data_im_in(31)=>mul_im_out(1013),
            data_im_in(32)=>mul_im_out(1045),
            data_im_in(33)=>mul_im_out(1077),
            data_im_in(34)=>mul_im_out(1109),
            data_im_in(35)=>mul_im_out(1141),
            data_im_in(36)=>mul_im_out(1173),
            data_im_in(37)=>mul_im_out(1205),
            data_im_in(38)=>mul_im_out(1237),
            data_im_in(39)=>mul_im_out(1269),
            data_im_in(40)=>mul_im_out(1301),
            data_im_in(41)=>mul_im_out(1333),
            data_im_in(42)=>mul_im_out(1365),
            data_im_in(43)=>mul_im_out(1397),
            data_im_in(44)=>mul_im_out(1429),
            data_im_in(45)=>mul_im_out(1461),
            data_im_in(46)=>mul_im_out(1493),
            data_im_in(47)=>mul_im_out(1525),
            data_im_in(48)=>mul_im_out(1557),
            data_im_in(49)=>mul_im_out(1589),
            data_im_in(50)=>mul_im_out(1621),
            data_im_in(51)=>mul_im_out(1653),
            data_im_in(52)=>mul_im_out(1685),
            data_im_in(53)=>mul_im_out(1717),
            data_im_in(54)=>mul_im_out(1749),
            data_im_in(55)=>mul_im_out(1781),
            data_im_in(56)=>mul_im_out(1813),
            data_im_in(57)=>mul_im_out(1845),
            data_im_in(58)=>mul_im_out(1877),
            data_im_in(59)=>mul_im_out(1909),
            data_im_in(60)=>mul_im_out(1941),
            data_im_in(61)=>mul_im_out(1973),
            data_im_in(62)=>mul_im_out(2005),
            data_im_in(63)=>mul_im_out(2037),
            data_re_out(0)=>data_re_out(21),
            data_re_out(1)=>data_re_out(53),
            data_re_out(2)=>data_re_out(85),
            data_re_out(3)=>data_re_out(117),
            data_re_out(4)=>data_re_out(149),
            data_re_out(5)=>data_re_out(181),
            data_re_out(6)=>data_re_out(213),
            data_re_out(7)=>data_re_out(245),
            data_re_out(8)=>data_re_out(277),
            data_re_out(9)=>data_re_out(309),
            data_re_out(10)=>data_re_out(341),
            data_re_out(11)=>data_re_out(373),
            data_re_out(12)=>data_re_out(405),
            data_re_out(13)=>data_re_out(437),
            data_re_out(14)=>data_re_out(469),
            data_re_out(15)=>data_re_out(501),
            data_re_out(16)=>data_re_out(533),
            data_re_out(17)=>data_re_out(565),
            data_re_out(18)=>data_re_out(597),
            data_re_out(19)=>data_re_out(629),
            data_re_out(20)=>data_re_out(661),
            data_re_out(21)=>data_re_out(693),
            data_re_out(22)=>data_re_out(725),
            data_re_out(23)=>data_re_out(757),
            data_re_out(24)=>data_re_out(789),
            data_re_out(25)=>data_re_out(821),
            data_re_out(26)=>data_re_out(853),
            data_re_out(27)=>data_re_out(885),
            data_re_out(28)=>data_re_out(917),
            data_re_out(29)=>data_re_out(949),
            data_re_out(30)=>data_re_out(981),
            data_re_out(31)=>data_re_out(1013),
            data_re_out(32)=>data_re_out(1045),
            data_re_out(33)=>data_re_out(1077),
            data_re_out(34)=>data_re_out(1109),
            data_re_out(35)=>data_re_out(1141),
            data_re_out(36)=>data_re_out(1173),
            data_re_out(37)=>data_re_out(1205),
            data_re_out(38)=>data_re_out(1237),
            data_re_out(39)=>data_re_out(1269),
            data_re_out(40)=>data_re_out(1301),
            data_re_out(41)=>data_re_out(1333),
            data_re_out(42)=>data_re_out(1365),
            data_re_out(43)=>data_re_out(1397),
            data_re_out(44)=>data_re_out(1429),
            data_re_out(45)=>data_re_out(1461),
            data_re_out(46)=>data_re_out(1493),
            data_re_out(47)=>data_re_out(1525),
            data_re_out(48)=>data_re_out(1557),
            data_re_out(49)=>data_re_out(1589),
            data_re_out(50)=>data_re_out(1621),
            data_re_out(51)=>data_re_out(1653),
            data_re_out(52)=>data_re_out(1685),
            data_re_out(53)=>data_re_out(1717),
            data_re_out(54)=>data_re_out(1749),
            data_re_out(55)=>data_re_out(1781),
            data_re_out(56)=>data_re_out(1813),
            data_re_out(57)=>data_re_out(1845),
            data_re_out(58)=>data_re_out(1877),
            data_re_out(59)=>data_re_out(1909),
            data_re_out(60)=>data_re_out(1941),
            data_re_out(61)=>data_re_out(1973),
            data_re_out(62)=>data_re_out(2005),
            data_re_out(63)=>data_re_out(2037),
            data_im_out(0)=>data_im_out(21),
            data_im_out(1)=>data_im_out(53),
            data_im_out(2)=>data_im_out(85),
            data_im_out(3)=>data_im_out(117),
            data_im_out(4)=>data_im_out(149),
            data_im_out(5)=>data_im_out(181),
            data_im_out(6)=>data_im_out(213),
            data_im_out(7)=>data_im_out(245),
            data_im_out(8)=>data_im_out(277),
            data_im_out(9)=>data_im_out(309),
            data_im_out(10)=>data_im_out(341),
            data_im_out(11)=>data_im_out(373),
            data_im_out(12)=>data_im_out(405),
            data_im_out(13)=>data_im_out(437),
            data_im_out(14)=>data_im_out(469),
            data_im_out(15)=>data_im_out(501),
            data_im_out(16)=>data_im_out(533),
            data_im_out(17)=>data_im_out(565),
            data_im_out(18)=>data_im_out(597),
            data_im_out(19)=>data_im_out(629),
            data_im_out(20)=>data_im_out(661),
            data_im_out(21)=>data_im_out(693),
            data_im_out(22)=>data_im_out(725),
            data_im_out(23)=>data_im_out(757),
            data_im_out(24)=>data_im_out(789),
            data_im_out(25)=>data_im_out(821),
            data_im_out(26)=>data_im_out(853),
            data_im_out(27)=>data_im_out(885),
            data_im_out(28)=>data_im_out(917),
            data_im_out(29)=>data_im_out(949),
            data_im_out(30)=>data_im_out(981),
            data_im_out(31)=>data_im_out(1013),
            data_im_out(32)=>data_im_out(1045),
            data_im_out(33)=>data_im_out(1077),
            data_im_out(34)=>data_im_out(1109),
            data_im_out(35)=>data_im_out(1141),
            data_im_out(36)=>data_im_out(1173),
            data_im_out(37)=>data_im_out(1205),
            data_im_out(38)=>data_im_out(1237),
            data_im_out(39)=>data_im_out(1269),
            data_im_out(40)=>data_im_out(1301),
            data_im_out(41)=>data_im_out(1333),
            data_im_out(42)=>data_im_out(1365),
            data_im_out(43)=>data_im_out(1397),
            data_im_out(44)=>data_im_out(1429),
            data_im_out(45)=>data_im_out(1461),
            data_im_out(46)=>data_im_out(1493),
            data_im_out(47)=>data_im_out(1525),
            data_im_out(48)=>data_im_out(1557),
            data_im_out(49)=>data_im_out(1589),
            data_im_out(50)=>data_im_out(1621),
            data_im_out(51)=>data_im_out(1653),
            data_im_out(52)=>data_im_out(1685),
            data_im_out(53)=>data_im_out(1717),
            data_im_out(54)=>data_im_out(1749),
            data_im_out(55)=>data_im_out(1781),
            data_im_out(56)=>data_im_out(1813),
            data_im_out(57)=>data_im_out(1845),
            data_im_out(58)=>data_im_out(1877),
            data_im_out(59)=>data_im_out(1909),
            data_im_out(60)=>data_im_out(1941),
            data_im_out(61)=>data_im_out(1973),
            data_im_out(62)=>data_im_out(2005),
            data_im_out(63)=>data_im_out(2037)
        );           

    URFFT_PT64_22 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(22),
            data_re_in(1)=>mul_re_out(54),
            data_re_in(2)=>mul_re_out(86),
            data_re_in(3)=>mul_re_out(118),
            data_re_in(4)=>mul_re_out(150),
            data_re_in(5)=>mul_re_out(182),
            data_re_in(6)=>mul_re_out(214),
            data_re_in(7)=>mul_re_out(246),
            data_re_in(8)=>mul_re_out(278),
            data_re_in(9)=>mul_re_out(310),
            data_re_in(10)=>mul_re_out(342),
            data_re_in(11)=>mul_re_out(374),
            data_re_in(12)=>mul_re_out(406),
            data_re_in(13)=>mul_re_out(438),
            data_re_in(14)=>mul_re_out(470),
            data_re_in(15)=>mul_re_out(502),
            data_re_in(16)=>mul_re_out(534),
            data_re_in(17)=>mul_re_out(566),
            data_re_in(18)=>mul_re_out(598),
            data_re_in(19)=>mul_re_out(630),
            data_re_in(20)=>mul_re_out(662),
            data_re_in(21)=>mul_re_out(694),
            data_re_in(22)=>mul_re_out(726),
            data_re_in(23)=>mul_re_out(758),
            data_re_in(24)=>mul_re_out(790),
            data_re_in(25)=>mul_re_out(822),
            data_re_in(26)=>mul_re_out(854),
            data_re_in(27)=>mul_re_out(886),
            data_re_in(28)=>mul_re_out(918),
            data_re_in(29)=>mul_re_out(950),
            data_re_in(30)=>mul_re_out(982),
            data_re_in(31)=>mul_re_out(1014),
            data_re_in(32)=>mul_re_out(1046),
            data_re_in(33)=>mul_re_out(1078),
            data_re_in(34)=>mul_re_out(1110),
            data_re_in(35)=>mul_re_out(1142),
            data_re_in(36)=>mul_re_out(1174),
            data_re_in(37)=>mul_re_out(1206),
            data_re_in(38)=>mul_re_out(1238),
            data_re_in(39)=>mul_re_out(1270),
            data_re_in(40)=>mul_re_out(1302),
            data_re_in(41)=>mul_re_out(1334),
            data_re_in(42)=>mul_re_out(1366),
            data_re_in(43)=>mul_re_out(1398),
            data_re_in(44)=>mul_re_out(1430),
            data_re_in(45)=>mul_re_out(1462),
            data_re_in(46)=>mul_re_out(1494),
            data_re_in(47)=>mul_re_out(1526),
            data_re_in(48)=>mul_re_out(1558),
            data_re_in(49)=>mul_re_out(1590),
            data_re_in(50)=>mul_re_out(1622),
            data_re_in(51)=>mul_re_out(1654),
            data_re_in(52)=>mul_re_out(1686),
            data_re_in(53)=>mul_re_out(1718),
            data_re_in(54)=>mul_re_out(1750),
            data_re_in(55)=>mul_re_out(1782),
            data_re_in(56)=>mul_re_out(1814),
            data_re_in(57)=>mul_re_out(1846),
            data_re_in(58)=>mul_re_out(1878),
            data_re_in(59)=>mul_re_out(1910),
            data_re_in(60)=>mul_re_out(1942),
            data_re_in(61)=>mul_re_out(1974),
            data_re_in(62)=>mul_re_out(2006),
            data_re_in(63)=>mul_re_out(2038),
            data_im_in(0)=>mul_im_out(22),
            data_im_in(1)=>mul_im_out(54),
            data_im_in(2)=>mul_im_out(86),
            data_im_in(3)=>mul_im_out(118),
            data_im_in(4)=>mul_im_out(150),
            data_im_in(5)=>mul_im_out(182),
            data_im_in(6)=>mul_im_out(214),
            data_im_in(7)=>mul_im_out(246),
            data_im_in(8)=>mul_im_out(278),
            data_im_in(9)=>mul_im_out(310),
            data_im_in(10)=>mul_im_out(342),
            data_im_in(11)=>mul_im_out(374),
            data_im_in(12)=>mul_im_out(406),
            data_im_in(13)=>mul_im_out(438),
            data_im_in(14)=>mul_im_out(470),
            data_im_in(15)=>mul_im_out(502),
            data_im_in(16)=>mul_im_out(534),
            data_im_in(17)=>mul_im_out(566),
            data_im_in(18)=>mul_im_out(598),
            data_im_in(19)=>mul_im_out(630),
            data_im_in(20)=>mul_im_out(662),
            data_im_in(21)=>mul_im_out(694),
            data_im_in(22)=>mul_im_out(726),
            data_im_in(23)=>mul_im_out(758),
            data_im_in(24)=>mul_im_out(790),
            data_im_in(25)=>mul_im_out(822),
            data_im_in(26)=>mul_im_out(854),
            data_im_in(27)=>mul_im_out(886),
            data_im_in(28)=>mul_im_out(918),
            data_im_in(29)=>mul_im_out(950),
            data_im_in(30)=>mul_im_out(982),
            data_im_in(31)=>mul_im_out(1014),
            data_im_in(32)=>mul_im_out(1046),
            data_im_in(33)=>mul_im_out(1078),
            data_im_in(34)=>mul_im_out(1110),
            data_im_in(35)=>mul_im_out(1142),
            data_im_in(36)=>mul_im_out(1174),
            data_im_in(37)=>mul_im_out(1206),
            data_im_in(38)=>mul_im_out(1238),
            data_im_in(39)=>mul_im_out(1270),
            data_im_in(40)=>mul_im_out(1302),
            data_im_in(41)=>mul_im_out(1334),
            data_im_in(42)=>mul_im_out(1366),
            data_im_in(43)=>mul_im_out(1398),
            data_im_in(44)=>mul_im_out(1430),
            data_im_in(45)=>mul_im_out(1462),
            data_im_in(46)=>mul_im_out(1494),
            data_im_in(47)=>mul_im_out(1526),
            data_im_in(48)=>mul_im_out(1558),
            data_im_in(49)=>mul_im_out(1590),
            data_im_in(50)=>mul_im_out(1622),
            data_im_in(51)=>mul_im_out(1654),
            data_im_in(52)=>mul_im_out(1686),
            data_im_in(53)=>mul_im_out(1718),
            data_im_in(54)=>mul_im_out(1750),
            data_im_in(55)=>mul_im_out(1782),
            data_im_in(56)=>mul_im_out(1814),
            data_im_in(57)=>mul_im_out(1846),
            data_im_in(58)=>mul_im_out(1878),
            data_im_in(59)=>mul_im_out(1910),
            data_im_in(60)=>mul_im_out(1942),
            data_im_in(61)=>mul_im_out(1974),
            data_im_in(62)=>mul_im_out(2006),
            data_im_in(63)=>mul_im_out(2038),
            data_re_out(0)=>data_re_out(22),
            data_re_out(1)=>data_re_out(54),
            data_re_out(2)=>data_re_out(86),
            data_re_out(3)=>data_re_out(118),
            data_re_out(4)=>data_re_out(150),
            data_re_out(5)=>data_re_out(182),
            data_re_out(6)=>data_re_out(214),
            data_re_out(7)=>data_re_out(246),
            data_re_out(8)=>data_re_out(278),
            data_re_out(9)=>data_re_out(310),
            data_re_out(10)=>data_re_out(342),
            data_re_out(11)=>data_re_out(374),
            data_re_out(12)=>data_re_out(406),
            data_re_out(13)=>data_re_out(438),
            data_re_out(14)=>data_re_out(470),
            data_re_out(15)=>data_re_out(502),
            data_re_out(16)=>data_re_out(534),
            data_re_out(17)=>data_re_out(566),
            data_re_out(18)=>data_re_out(598),
            data_re_out(19)=>data_re_out(630),
            data_re_out(20)=>data_re_out(662),
            data_re_out(21)=>data_re_out(694),
            data_re_out(22)=>data_re_out(726),
            data_re_out(23)=>data_re_out(758),
            data_re_out(24)=>data_re_out(790),
            data_re_out(25)=>data_re_out(822),
            data_re_out(26)=>data_re_out(854),
            data_re_out(27)=>data_re_out(886),
            data_re_out(28)=>data_re_out(918),
            data_re_out(29)=>data_re_out(950),
            data_re_out(30)=>data_re_out(982),
            data_re_out(31)=>data_re_out(1014),
            data_re_out(32)=>data_re_out(1046),
            data_re_out(33)=>data_re_out(1078),
            data_re_out(34)=>data_re_out(1110),
            data_re_out(35)=>data_re_out(1142),
            data_re_out(36)=>data_re_out(1174),
            data_re_out(37)=>data_re_out(1206),
            data_re_out(38)=>data_re_out(1238),
            data_re_out(39)=>data_re_out(1270),
            data_re_out(40)=>data_re_out(1302),
            data_re_out(41)=>data_re_out(1334),
            data_re_out(42)=>data_re_out(1366),
            data_re_out(43)=>data_re_out(1398),
            data_re_out(44)=>data_re_out(1430),
            data_re_out(45)=>data_re_out(1462),
            data_re_out(46)=>data_re_out(1494),
            data_re_out(47)=>data_re_out(1526),
            data_re_out(48)=>data_re_out(1558),
            data_re_out(49)=>data_re_out(1590),
            data_re_out(50)=>data_re_out(1622),
            data_re_out(51)=>data_re_out(1654),
            data_re_out(52)=>data_re_out(1686),
            data_re_out(53)=>data_re_out(1718),
            data_re_out(54)=>data_re_out(1750),
            data_re_out(55)=>data_re_out(1782),
            data_re_out(56)=>data_re_out(1814),
            data_re_out(57)=>data_re_out(1846),
            data_re_out(58)=>data_re_out(1878),
            data_re_out(59)=>data_re_out(1910),
            data_re_out(60)=>data_re_out(1942),
            data_re_out(61)=>data_re_out(1974),
            data_re_out(62)=>data_re_out(2006),
            data_re_out(63)=>data_re_out(2038),
            data_im_out(0)=>data_im_out(22),
            data_im_out(1)=>data_im_out(54),
            data_im_out(2)=>data_im_out(86),
            data_im_out(3)=>data_im_out(118),
            data_im_out(4)=>data_im_out(150),
            data_im_out(5)=>data_im_out(182),
            data_im_out(6)=>data_im_out(214),
            data_im_out(7)=>data_im_out(246),
            data_im_out(8)=>data_im_out(278),
            data_im_out(9)=>data_im_out(310),
            data_im_out(10)=>data_im_out(342),
            data_im_out(11)=>data_im_out(374),
            data_im_out(12)=>data_im_out(406),
            data_im_out(13)=>data_im_out(438),
            data_im_out(14)=>data_im_out(470),
            data_im_out(15)=>data_im_out(502),
            data_im_out(16)=>data_im_out(534),
            data_im_out(17)=>data_im_out(566),
            data_im_out(18)=>data_im_out(598),
            data_im_out(19)=>data_im_out(630),
            data_im_out(20)=>data_im_out(662),
            data_im_out(21)=>data_im_out(694),
            data_im_out(22)=>data_im_out(726),
            data_im_out(23)=>data_im_out(758),
            data_im_out(24)=>data_im_out(790),
            data_im_out(25)=>data_im_out(822),
            data_im_out(26)=>data_im_out(854),
            data_im_out(27)=>data_im_out(886),
            data_im_out(28)=>data_im_out(918),
            data_im_out(29)=>data_im_out(950),
            data_im_out(30)=>data_im_out(982),
            data_im_out(31)=>data_im_out(1014),
            data_im_out(32)=>data_im_out(1046),
            data_im_out(33)=>data_im_out(1078),
            data_im_out(34)=>data_im_out(1110),
            data_im_out(35)=>data_im_out(1142),
            data_im_out(36)=>data_im_out(1174),
            data_im_out(37)=>data_im_out(1206),
            data_im_out(38)=>data_im_out(1238),
            data_im_out(39)=>data_im_out(1270),
            data_im_out(40)=>data_im_out(1302),
            data_im_out(41)=>data_im_out(1334),
            data_im_out(42)=>data_im_out(1366),
            data_im_out(43)=>data_im_out(1398),
            data_im_out(44)=>data_im_out(1430),
            data_im_out(45)=>data_im_out(1462),
            data_im_out(46)=>data_im_out(1494),
            data_im_out(47)=>data_im_out(1526),
            data_im_out(48)=>data_im_out(1558),
            data_im_out(49)=>data_im_out(1590),
            data_im_out(50)=>data_im_out(1622),
            data_im_out(51)=>data_im_out(1654),
            data_im_out(52)=>data_im_out(1686),
            data_im_out(53)=>data_im_out(1718),
            data_im_out(54)=>data_im_out(1750),
            data_im_out(55)=>data_im_out(1782),
            data_im_out(56)=>data_im_out(1814),
            data_im_out(57)=>data_im_out(1846),
            data_im_out(58)=>data_im_out(1878),
            data_im_out(59)=>data_im_out(1910),
            data_im_out(60)=>data_im_out(1942),
            data_im_out(61)=>data_im_out(1974),
            data_im_out(62)=>data_im_out(2006),
            data_im_out(63)=>data_im_out(2038)
        );           

    URFFT_PT64_23 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(23),
            data_re_in(1)=>mul_re_out(55),
            data_re_in(2)=>mul_re_out(87),
            data_re_in(3)=>mul_re_out(119),
            data_re_in(4)=>mul_re_out(151),
            data_re_in(5)=>mul_re_out(183),
            data_re_in(6)=>mul_re_out(215),
            data_re_in(7)=>mul_re_out(247),
            data_re_in(8)=>mul_re_out(279),
            data_re_in(9)=>mul_re_out(311),
            data_re_in(10)=>mul_re_out(343),
            data_re_in(11)=>mul_re_out(375),
            data_re_in(12)=>mul_re_out(407),
            data_re_in(13)=>mul_re_out(439),
            data_re_in(14)=>mul_re_out(471),
            data_re_in(15)=>mul_re_out(503),
            data_re_in(16)=>mul_re_out(535),
            data_re_in(17)=>mul_re_out(567),
            data_re_in(18)=>mul_re_out(599),
            data_re_in(19)=>mul_re_out(631),
            data_re_in(20)=>mul_re_out(663),
            data_re_in(21)=>mul_re_out(695),
            data_re_in(22)=>mul_re_out(727),
            data_re_in(23)=>mul_re_out(759),
            data_re_in(24)=>mul_re_out(791),
            data_re_in(25)=>mul_re_out(823),
            data_re_in(26)=>mul_re_out(855),
            data_re_in(27)=>mul_re_out(887),
            data_re_in(28)=>mul_re_out(919),
            data_re_in(29)=>mul_re_out(951),
            data_re_in(30)=>mul_re_out(983),
            data_re_in(31)=>mul_re_out(1015),
            data_re_in(32)=>mul_re_out(1047),
            data_re_in(33)=>mul_re_out(1079),
            data_re_in(34)=>mul_re_out(1111),
            data_re_in(35)=>mul_re_out(1143),
            data_re_in(36)=>mul_re_out(1175),
            data_re_in(37)=>mul_re_out(1207),
            data_re_in(38)=>mul_re_out(1239),
            data_re_in(39)=>mul_re_out(1271),
            data_re_in(40)=>mul_re_out(1303),
            data_re_in(41)=>mul_re_out(1335),
            data_re_in(42)=>mul_re_out(1367),
            data_re_in(43)=>mul_re_out(1399),
            data_re_in(44)=>mul_re_out(1431),
            data_re_in(45)=>mul_re_out(1463),
            data_re_in(46)=>mul_re_out(1495),
            data_re_in(47)=>mul_re_out(1527),
            data_re_in(48)=>mul_re_out(1559),
            data_re_in(49)=>mul_re_out(1591),
            data_re_in(50)=>mul_re_out(1623),
            data_re_in(51)=>mul_re_out(1655),
            data_re_in(52)=>mul_re_out(1687),
            data_re_in(53)=>mul_re_out(1719),
            data_re_in(54)=>mul_re_out(1751),
            data_re_in(55)=>mul_re_out(1783),
            data_re_in(56)=>mul_re_out(1815),
            data_re_in(57)=>mul_re_out(1847),
            data_re_in(58)=>mul_re_out(1879),
            data_re_in(59)=>mul_re_out(1911),
            data_re_in(60)=>mul_re_out(1943),
            data_re_in(61)=>mul_re_out(1975),
            data_re_in(62)=>mul_re_out(2007),
            data_re_in(63)=>mul_re_out(2039),
            data_im_in(0)=>mul_im_out(23),
            data_im_in(1)=>mul_im_out(55),
            data_im_in(2)=>mul_im_out(87),
            data_im_in(3)=>mul_im_out(119),
            data_im_in(4)=>mul_im_out(151),
            data_im_in(5)=>mul_im_out(183),
            data_im_in(6)=>mul_im_out(215),
            data_im_in(7)=>mul_im_out(247),
            data_im_in(8)=>mul_im_out(279),
            data_im_in(9)=>mul_im_out(311),
            data_im_in(10)=>mul_im_out(343),
            data_im_in(11)=>mul_im_out(375),
            data_im_in(12)=>mul_im_out(407),
            data_im_in(13)=>mul_im_out(439),
            data_im_in(14)=>mul_im_out(471),
            data_im_in(15)=>mul_im_out(503),
            data_im_in(16)=>mul_im_out(535),
            data_im_in(17)=>mul_im_out(567),
            data_im_in(18)=>mul_im_out(599),
            data_im_in(19)=>mul_im_out(631),
            data_im_in(20)=>mul_im_out(663),
            data_im_in(21)=>mul_im_out(695),
            data_im_in(22)=>mul_im_out(727),
            data_im_in(23)=>mul_im_out(759),
            data_im_in(24)=>mul_im_out(791),
            data_im_in(25)=>mul_im_out(823),
            data_im_in(26)=>mul_im_out(855),
            data_im_in(27)=>mul_im_out(887),
            data_im_in(28)=>mul_im_out(919),
            data_im_in(29)=>mul_im_out(951),
            data_im_in(30)=>mul_im_out(983),
            data_im_in(31)=>mul_im_out(1015),
            data_im_in(32)=>mul_im_out(1047),
            data_im_in(33)=>mul_im_out(1079),
            data_im_in(34)=>mul_im_out(1111),
            data_im_in(35)=>mul_im_out(1143),
            data_im_in(36)=>mul_im_out(1175),
            data_im_in(37)=>mul_im_out(1207),
            data_im_in(38)=>mul_im_out(1239),
            data_im_in(39)=>mul_im_out(1271),
            data_im_in(40)=>mul_im_out(1303),
            data_im_in(41)=>mul_im_out(1335),
            data_im_in(42)=>mul_im_out(1367),
            data_im_in(43)=>mul_im_out(1399),
            data_im_in(44)=>mul_im_out(1431),
            data_im_in(45)=>mul_im_out(1463),
            data_im_in(46)=>mul_im_out(1495),
            data_im_in(47)=>mul_im_out(1527),
            data_im_in(48)=>mul_im_out(1559),
            data_im_in(49)=>mul_im_out(1591),
            data_im_in(50)=>mul_im_out(1623),
            data_im_in(51)=>mul_im_out(1655),
            data_im_in(52)=>mul_im_out(1687),
            data_im_in(53)=>mul_im_out(1719),
            data_im_in(54)=>mul_im_out(1751),
            data_im_in(55)=>mul_im_out(1783),
            data_im_in(56)=>mul_im_out(1815),
            data_im_in(57)=>mul_im_out(1847),
            data_im_in(58)=>mul_im_out(1879),
            data_im_in(59)=>mul_im_out(1911),
            data_im_in(60)=>mul_im_out(1943),
            data_im_in(61)=>mul_im_out(1975),
            data_im_in(62)=>mul_im_out(2007),
            data_im_in(63)=>mul_im_out(2039),
            data_re_out(0)=>data_re_out(23),
            data_re_out(1)=>data_re_out(55),
            data_re_out(2)=>data_re_out(87),
            data_re_out(3)=>data_re_out(119),
            data_re_out(4)=>data_re_out(151),
            data_re_out(5)=>data_re_out(183),
            data_re_out(6)=>data_re_out(215),
            data_re_out(7)=>data_re_out(247),
            data_re_out(8)=>data_re_out(279),
            data_re_out(9)=>data_re_out(311),
            data_re_out(10)=>data_re_out(343),
            data_re_out(11)=>data_re_out(375),
            data_re_out(12)=>data_re_out(407),
            data_re_out(13)=>data_re_out(439),
            data_re_out(14)=>data_re_out(471),
            data_re_out(15)=>data_re_out(503),
            data_re_out(16)=>data_re_out(535),
            data_re_out(17)=>data_re_out(567),
            data_re_out(18)=>data_re_out(599),
            data_re_out(19)=>data_re_out(631),
            data_re_out(20)=>data_re_out(663),
            data_re_out(21)=>data_re_out(695),
            data_re_out(22)=>data_re_out(727),
            data_re_out(23)=>data_re_out(759),
            data_re_out(24)=>data_re_out(791),
            data_re_out(25)=>data_re_out(823),
            data_re_out(26)=>data_re_out(855),
            data_re_out(27)=>data_re_out(887),
            data_re_out(28)=>data_re_out(919),
            data_re_out(29)=>data_re_out(951),
            data_re_out(30)=>data_re_out(983),
            data_re_out(31)=>data_re_out(1015),
            data_re_out(32)=>data_re_out(1047),
            data_re_out(33)=>data_re_out(1079),
            data_re_out(34)=>data_re_out(1111),
            data_re_out(35)=>data_re_out(1143),
            data_re_out(36)=>data_re_out(1175),
            data_re_out(37)=>data_re_out(1207),
            data_re_out(38)=>data_re_out(1239),
            data_re_out(39)=>data_re_out(1271),
            data_re_out(40)=>data_re_out(1303),
            data_re_out(41)=>data_re_out(1335),
            data_re_out(42)=>data_re_out(1367),
            data_re_out(43)=>data_re_out(1399),
            data_re_out(44)=>data_re_out(1431),
            data_re_out(45)=>data_re_out(1463),
            data_re_out(46)=>data_re_out(1495),
            data_re_out(47)=>data_re_out(1527),
            data_re_out(48)=>data_re_out(1559),
            data_re_out(49)=>data_re_out(1591),
            data_re_out(50)=>data_re_out(1623),
            data_re_out(51)=>data_re_out(1655),
            data_re_out(52)=>data_re_out(1687),
            data_re_out(53)=>data_re_out(1719),
            data_re_out(54)=>data_re_out(1751),
            data_re_out(55)=>data_re_out(1783),
            data_re_out(56)=>data_re_out(1815),
            data_re_out(57)=>data_re_out(1847),
            data_re_out(58)=>data_re_out(1879),
            data_re_out(59)=>data_re_out(1911),
            data_re_out(60)=>data_re_out(1943),
            data_re_out(61)=>data_re_out(1975),
            data_re_out(62)=>data_re_out(2007),
            data_re_out(63)=>data_re_out(2039),
            data_im_out(0)=>data_im_out(23),
            data_im_out(1)=>data_im_out(55),
            data_im_out(2)=>data_im_out(87),
            data_im_out(3)=>data_im_out(119),
            data_im_out(4)=>data_im_out(151),
            data_im_out(5)=>data_im_out(183),
            data_im_out(6)=>data_im_out(215),
            data_im_out(7)=>data_im_out(247),
            data_im_out(8)=>data_im_out(279),
            data_im_out(9)=>data_im_out(311),
            data_im_out(10)=>data_im_out(343),
            data_im_out(11)=>data_im_out(375),
            data_im_out(12)=>data_im_out(407),
            data_im_out(13)=>data_im_out(439),
            data_im_out(14)=>data_im_out(471),
            data_im_out(15)=>data_im_out(503),
            data_im_out(16)=>data_im_out(535),
            data_im_out(17)=>data_im_out(567),
            data_im_out(18)=>data_im_out(599),
            data_im_out(19)=>data_im_out(631),
            data_im_out(20)=>data_im_out(663),
            data_im_out(21)=>data_im_out(695),
            data_im_out(22)=>data_im_out(727),
            data_im_out(23)=>data_im_out(759),
            data_im_out(24)=>data_im_out(791),
            data_im_out(25)=>data_im_out(823),
            data_im_out(26)=>data_im_out(855),
            data_im_out(27)=>data_im_out(887),
            data_im_out(28)=>data_im_out(919),
            data_im_out(29)=>data_im_out(951),
            data_im_out(30)=>data_im_out(983),
            data_im_out(31)=>data_im_out(1015),
            data_im_out(32)=>data_im_out(1047),
            data_im_out(33)=>data_im_out(1079),
            data_im_out(34)=>data_im_out(1111),
            data_im_out(35)=>data_im_out(1143),
            data_im_out(36)=>data_im_out(1175),
            data_im_out(37)=>data_im_out(1207),
            data_im_out(38)=>data_im_out(1239),
            data_im_out(39)=>data_im_out(1271),
            data_im_out(40)=>data_im_out(1303),
            data_im_out(41)=>data_im_out(1335),
            data_im_out(42)=>data_im_out(1367),
            data_im_out(43)=>data_im_out(1399),
            data_im_out(44)=>data_im_out(1431),
            data_im_out(45)=>data_im_out(1463),
            data_im_out(46)=>data_im_out(1495),
            data_im_out(47)=>data_im_out(1527),
            data_im_out(48)=>data_im_out(1559),
            data_im_out(49)=>data_im_out(1591),
            data_im_out(50)=>data_im_out(1623),
            data_im_out(51)=>data_im_out(1655),
            data_im_out(52)=>data_im_out(1687),
            data_im_out(53)=>data_im_out(1719),
            data_im_out(54)=>data_im_out(1751),
            data_im_out(55)=>data_im_out(1783),
            data_im_out(56)=>data_im_out(1815),
            data_im_out(57)=>data_im_out(1847),
            data_im_out(58)=>data_im_out(1879),
            data_im_out(59)=>data_im_out(1911),
            data_im_out(60)=>data_im_out(1943),
            data_im_out(61)=>data_im_out(1975),
            data_im_out(62)=>data_im_out(2007),
            data_im_out(63)=>data_im_out(2039)
        );           

    URFFT_PT64_24 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(24),
            data_re_in(1)=>mul_re_out(56),
            data_re_in(2)=>mul_re_out(88),
            data_re_in(3)=>mul_re_out(120),
            data_re_in(4)=>mul_re_out(152),
            data_re_in(5)=>mul_re_out(184),
            data_re_in(6)=>mul_re_out(216),
            data_re_in(7)=>mul_re_out(248),
            data_re_in(8)=>mul_re_out(280),
            data_re_in(9)=>mul_re_out(312),
            data_re_in(10)=>mul_re_out(344),
            data_re_in(11)=>mul_re_out(376),
            data_re_in(12)=>mul_re_out(408),
            data_re_in(13)=>mul_re_out(440),
            data_re_in(14)=>mul_re_out(472),
            data_re_in(15)=>mul_re_out(504),
            data_re_in(16)=>mul_re_out(536),
            data_re_in(17)=>mul_re_out(568),
            data_re_in(18)=>mul_re_out(600),
            data_re_in(19)=>mul_re_out(632),
            data_re_in(20)=>mul_re_out(664),
            data_re_in(21)=>mul_re_out(696),
            data_re_in(22)=>mul_re_out(728),
            data_re_in(23)=>mul_re_out(760),
            data_re_in(24)=>mul_re_out(792),
            data_re_in(25)=>mul_re_out(824),
            data_re_in(26)=>mul_re_out(856),
            data_re_in(27)=>mul_re_out(888),
            data_re_in(28)=>mul_re_out(920),
            data_re_in(29)=>mul_re_out(952),
            data_re_in(30)=>mul_re_out(984),
            data_re_in(31)=>mul_re_out(1016),
            data_re_in(32)=>mul_re_out(1048),
            data_re_in(33)=>mul_re_out(1080),
            data_re_in(34)=>mul_re_out(1112),
            data_re_in(35)=>mul_re_out(1144),
            data_re_in(36)=>mul_re_out(1176),
            data_re_in(37)=>mul_re_out(1208),
            data_re_in(38)=>mul_re_out(1240),
            data_re_in(39)=>mul_re_out(1272),
            data_re_in(40)=>mul_re_out(1304),
            data_re_in(41)=>mul_re_out(1336),
            data_re_in(42)=>mul_re_out(1368),
            data_re_in(43)=>mul_re_out(1400),
            data_re_in(44)=>mul_re_out(1432),
            data_re_in(45)=>mul_re_out(1464),
            data_re_in(46)=>mul_re_out(1496),
            data_re_in(47)=>mul_re_out(1528),
            data_re_in(48)=>mul_re_out(1560),
            data_re_in(49)=>mul_re_out(1592),
            data_re_in(50)=>mul_re_out(1624),
            data_re_in(51)=>mul_re_out(1656),
            data_re_in(52)=>mul_re_out(1688),
            data_re_in(53)=>mul_re_out(1720),
            data_re_in(54)=>mul_re_out(1752),
            data_re_in(55)=>mul_re_out(1784),
            data_re_in(56)=>mul_re_out(1816),
            data_re_in(57)=>mul_re_out(1848),
            data_re_in(58)=>mul_re_out(1880),
            data_re_in(59)=>mul_re_out(1912),
            data_re_in(60)=>mul_re_out(1944),
            data_re_in(61)=>mul_re_out(1976),
            data_re_in(62)=>mul_re_out(2008),
            data_re_in(63)=>mul_re_out(2040),
            data_im_in(0)=>mul_im_out(24),
            data_im_in(1)=>mul_im_out(56),
            data_im_in(2)=>mul_im_out(88),
            data_im_in(3)=>mul_im_out(120),
            data_im_in(4)=>mul_im_out(152),
            data_im_in(5)=>mul_im_out(184),
            data_im_in(6)=>mul_im_out(216),
            data_im_in(7)=>mul_im_out(248),
            data_im_in(8)=>mul_im_out(280),
            data_im_in(9)=>mul_im_out(312),
            data_im_in(10)=>mul_im_out(344),
            data_im_in(11)=>mul_im_out(376),
            data_im_in(12)=>mul_im_out(408),
            data_im_in(13)=>mul_im_out(440),
            data_im_in(14)=>mul_im_out(472),
            data_im_in(15)=>mul_im_out(504),
            data_im_in(16)=>mul_im_out(536),
            data_im_in(17)=>mul_im_out(568),
            data_im_in(18)=>mul_im_out(600),
            data_im_in(19)=>mul_im_out(632),
            data_im_in(20)=>mul_im_out(664),
            data_im_in(21)=>mul_im_out(696),
            data_im_in(22)=>mul_im_out(728),
            data_im_in(23)=>mul_im_out(760),
            data_im_in(24)=>mul_im_out(792),
            data_im_in(25)=>mul_im_out(824),
            data_im_in(26)=>mul_im_out(856),
            data_im_in(27)=>mul_im_out(888),
            data_im_in(28)=>mul_im_out(920),
            data_im_in(29)=>mul_im_out(952),
            data_im_in(30)=>mul_im_out(984),
            data_im_in(31)=>mul_im_out(1016),
            data_im_in(32)=>mul_im_out(1048),
            data_im_in(33)=>mul_im_out(1080),
            data_im_in(34)=>mul_im_out(1112),
            data_im_in(35)=>mul_im_out(1144),
            data_im_in(36)=>mul_im_out(1176),
            data_im_in(37)=>mul_im_out(1208),
            data_im_in(38)=>mul_im_out(1240),
            data_im_in(39)=>mul_im_out(1272),
            data_im_in(40)=>mul_im_out(1304),
            data_im_in(41)=>mul_im_out(1336),
            data_im_in(42)=>mul_im_out(1368),
            data_im_in(43)=>mul_im_out(1400),
            data_im_in(44)=>mul_im_out(1432),
            data_im_in(45)=>mul_im_out(1464),
            data_im_in(46)=>mul_im_out(1496),
            data_im_in(47)=>mul_im_out(1528),
            data_im_in(48)=>mul_im_out(1560),
            data_im_in(49)=>mul_im_out(1592),
            data_im_in(50)=>mul_im_out(1624),
            data_im_in(51)=>mul_im_out(1656),
            data_im_in(52)=>mul_im_out(1688),
            data_im_in(53)=>mul_im_out(1720),
            data_im_in(54)=>mul_im_out(1752),
            data_im_in(55)=>mul_im_out(1784),
            data_im_in(56)=>mul_im_out(1816),
            data_im_in(57)=>mul_im_out(1848),
            data_im_in(58)=>mul_im_out(1880),
            data_im_in(59)=>mul_im_out(1912),
            data_im_in(60)=>mul_im_out(1944),
            data_im_in(61)=>mul_im_out(1976),
            data_im_in(62)=>mul_im_out(2008),
            data_im_in(63)=>mul_im_out(2040),
            data_re_out(0)=>data_re_out(24),
            data_re_out(1)=>data_re_out(56),
            data_re_out(2)=>data_re_out(88),
            data_re_out(3)=>data_re_out(120),
            data_re_out(4)=>data_re_out(152),
            data_re_out(5)=>data_re_out(184),
            data_re_out(6)=>data_re_out(216),
            data_re_out(7)=>data_re_out(248),
            data_re_out(8)=>data_re_out(280),
            data_re_out(9)=>data_re_out(312),
            data_re_out(10)=>data_re_out(344),
            data_re_out(11)=>data_re_out(376),
            data_re_out(12)=>data_re_out(408),
            data_re_out(13)=>data_re_out(440),
            data_re_out(14)=>data_re_out(472),
            data_re_out(15)=>data_re_out(504),
            data_re_out(16)=>data_re_out(536),
            data_re_out(17)=>data_re_out(568),
            data_re_out(18)=>data_re_out(600),
            data_re_out(19)=>data_re_out(632),
            data_re_out(20)=>data_re_out(664),
            data_re_out(21)=>data_re_out(696),
            data_re_out(22)=>data_re_out(728),
            data_re_out(23)=>data_re_out(760),
            data_re_out(24)=>data_re_out(792),
            data_re_out(25)=>data_re_out(824),
            data_re_out(26)=>data_re_out(856),
            data_re_out(27)=>data_re_out(888),
            data_re_out(28)=>data_re_out(920),
            data_re_out(29)=>data_re_out(952),
            data_re_out(30)=>data_re_out(984),
            data_re_out(31)=>data_re_out(1016),
            data_re_out(32)=>data_re_out(1048),
            data_re_out(33)=>data_re_out(1080),
            data_re_out(34)=>data_re_out(1112),
            data_re_out(35)=>data_re_out(1144),
            data_re_out(36)=>data_re_out(1176),
            data_re_out(37)=>data_re_out(1208),
            data_re_out(38)=>data_re_out(1240),
            data_re_out(39)=>data_re_out(1272),
            data_re_out(40)=>data_re_out(1304),
            data_re_out(41)=>data_re_out(1336),
            data_re_out(42)=>data_re_out(1368),
            data_re_out(43)=>data_re_out(1400),
            data_re_out(44)=>data_re_out(1432),
            data_re_out(45)=>data_re_out(1464),
            data_re_out(46)=>data_re_out(1496),
            data_re_out(47)=>data_re_out(1528),
            data_re_out(48)=>data_re_out(1560),
            data_re_out(49)=>data_re_out(1592),
            data_re_out(50)=>data_re_out(1624),
            data_re_out(51)=>data_re_out(1656),
            data_re_out(52)=>data_re_out(1688),
            data_re_out(53)=>data_re_out(1720),
            data_re_out(54)=>data_re_out(1752),
            data_re_out(55)=>data_re_out(1784),
            data_re_out(56)=>data_re_out(1816),
            data_re_out(57)=>data_re_out(1848),
            data_re_out(58)=>data_re_out(1880),
            data_re_out(59)=>data_re_out(1912),
            data_re_out(60)=>data_re_out(1944),
            data_re_out(61)=>data_re_out(1976),
            data_re_out(62)=>data_re_out(2008),
            data_re_out(63)=>data_re_out(2040),
            data_im_out(0)=>data_im_out(24),
            data_im_out(1)=>data_im_out(56),
            data_im_out(2)=>data_im_out(88),
            data_im_out(3)=>data_im_out(120),
            data_im_out(4)=>data_im_out(152),
            data_im_out(5)=>data_im_out(184),
            data_im_out(6)=>data_im_out(216),
            data_im_out(7)=>data_im_out(248),
            data_im_out(8)=>data_im_out(280),
            data_im_out(9)=>data_im_out(312),
            data_im_out(10)=>data_im_out(344),
            data_im_out(11)=>data_im_out(376),
            data_im_out(12)=>data_im_out(408),
            data_im_out(13)=>data_im_out(440),
            data_im_out(14)=>data_im_out(472),
            data_im_out(15)=>data_im_out(504),
            data_im_out(16)=>data_im_out(536),
            data_im_out(17)=>data_im_out(568),
            data_im_out(18)=>data_im_out(600),
            data_im_out(19)=>data_im_out(632),
            data_im_out(20)=>data_im_out(664),
            data_im_out(21)=>data_im_out(696),
            data_im_out(22)=>data_im_out(728),
            data_im_out(23)=>data_im_out(760),
            data_im_out(24)=>data_im_out(792),
            data_im_out(25)=>data_im_out(824),
            data_im_out(26)=>data_im_out(856),
            data_im_out(27)=>data_im_out(888),
            data_im_out(28)=>data_im_out(920),
            data_im_out(29)=>data_im_out(952),
            data_im_out(30)=>data_im_out(984),
            data_im_out(31)=>data_im_out(1016),
            data_im_out(32)=>data_im_out(1048),
            data_im_out(33)=>data_im_out(1080),
            data_im_out(34)=>data_im_out(1112),
            data_im_out(35)=>data_im_out(1144),
            data_im_out(36)=>data_im_out(1176),
            data_im_out(37)=>data_im_out(1208),
            data_im_out(38)=>data_im_out(1240),
            data_im_out(39)=>data_im_out(1272),
            data_im_out(40)=>data_im_out(1304),
            data_im_out(41)=>data_im_out(1336),
            data_im_out(42)=>data_im_out(1368),
            data_im_out(43)=>data_im_out(1400),
            data_im_out(44)=>data_im_out(1432),
            data_im_out(45)=>data_im_out(1464),
            data_im_out(46)=>data_im_out(1496),
            data_im_out(47)=>data_im_out(1528),
            data_im_out(48)=>data_im_out(1560),
            data_im_out(49)=>data_im_out(1592),
            data_im_out(50)=>data_im_out(1624),
            data_im_out(51)=>data_im_out(1656),
            data_im_out(52)=>data_im_out(1688),
            data_im_out(53)=>data_im_out(1720),
            data_im_out(54)=>data_im_out(1752),
            data_im_out(55)=>data_im_out(1784),
            data_im_out(56)=>data_im_out(1816),
            data_im_out(57)=>data_im_out(1848),
            data_im_out(58)=>data_im_out(1880),
            data_im_out(59)=>data_im_out(1912),
            data_im_out(60)=>data_im_out(1944),
            data_im_out(61)=>data_im_out(1976),
            data_im_out(62)=>data_im_out(2008),
            data_im_out(63)=>data_im_out(2040)
        );           

    URFFT_PT64_25 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(25),
            data_re_in(1)=>mul_re_out(57),
            data_re_in(2)=>mul_re_out(89),
            data_re_in(3)=>mul_re_out(121),
            data_re_in(4)=>mul_re_out(153),
            data_re_in(5)=>mul_re_out(185),
            data_re_in(6)=>mul_re_out(217),
            data_re_in(7)=>mul_re_out(249),
            data_re_in(8)=>mul_re_out(281),
            data_re_in(9)=>mul_re_out(313),
            data_re_in(10)=>mul_re_out(345),
            data_re_in(11)=>mul_re_out(377),
            data_re_in(12)=>mul_re_out(409),
            data_re_in(13)=>mul_re_out(441),
            data_re_in(14)=>mul_re_out(473),
            data_re_in(15)=>mul_re_out(505),
            data_re_in(16)=>mul_re_out(537),
            data_re_in(17)=>mul_re_out(569),
            data_re_in(18)=>mul_re_out(601),
            data_re_in(19)=>mul_re_out(633),
            data_re_in(20)=>mul_re_out(665),
            data_re_in(21)=>mul_re_out(697),
            data_re_in(22)=>mul_re_out(729),
            data_re_in(23)=>mul_re_out(761),
            data_re_in(24)=>mul_re_out(793),
            data_re_in(25)=>mul_re_out(825),
            data_re_in(26)=>mul_re_out(857),
            data_re_in(27)=>mul_re_out(889),
            data_re_in(28)=>mul_re_out(921),
            data_re_in(29)=>mul_re_out(953),
            data_re_in(30)=>mul_re_out(985),
            data_re_in(31)=>mul_re_out(1017),
            data_re_in(32)=>mul_re_out(1049),
            data_re_in(33)=>mul_re_out(1081),
            data_re_in(34)=>mul_re_out(1113),
            data_re_in(35)=>mul_re_out(1145),
            data_re_in(36)=>mul_re_out(1177),
            data_re_in(37)=>mul_re_out(1209),
            data_re_in(38)=>mul_re_out(1241),
            data_re_in(39)=>mul_re_out(1273),
            data_re_in(40)=>mul_re_out(1305),
            data_re_in(41)=>mul_re_out(1337),
            data_re_in(42)=>mul_re_out(1369),
            data_re_in(43)=>mul_re_out(1401),
            data_re_in(44)=>mul_re_out(1433),
            data_re_in(45)=>mul_re_out(1465),
            data_re_in(46)=>mul_re_out(1497),
            data_re_in(47)=>mul_re_out(1529),
            data_re_in(48)=>mul_re_out(1561),
            data_re_in(49)=>mul_re_out(1593),
            data_re_in(50)=>mul_re_out(1625),
            data_re_in(51)=>mul_re_out(1657),
            data_re_in(52)=>mul_re_out(1689),
            data_re_in(53)=>mul_re_out(1721),
            data_re_in(54)=>mul_re_out(1753),
            data_re_in(55)=>mul_re_out(1785),
            data_re_in(56)=>mul_re_out(1817),
            data_re_in(57)=>mul_re_out(1849),
            data_re_in(58)=>mul_re_out(1881),
            data_re_in(59)=>mul_re_out(1913),
            data_re_in(60)=>mul_re_out(1945),
            data_re_in(61)=>mul_re_out(1977),
            data_re_in(62)=>mul_re_out(2009),
            data_re_in(63)=>mul_re_out(2041),
            data_im_in(0)=>mul_im_out(25),
            data_im_in(1)=>mul_im_out(57),
            data_im_in(2)=>mul_im_out(89),
            data_im_in(3)=>mul_im_out(121),
            data_im_in(4)=>mul_im_out(153),
            data_im_in(5)=>mul_im_out(185),
            data_im_in(6)=>mul_im_out(217),
            data_im_in(7)=>mul_im_out(249),
            data_im_in(8)=>mul_im_out(281),
            data_im_in(9)=>mul_im_out(313),
            data_im_in(10)=>mul_im_out(345),
            data_im_in(11)=>mul_im_out(377),
            data_im_in(12)=>mul_im_out(409),
            data_im_in(13)=>mul_im_out(441),
            data_im_in(14)=>mul_im_out(473),
            data_im_in(15)=>mul_im_out(505),
            data_im_in(16)=>mul_im_out(537),
            data_im_in(17)=>mul_im_out(569),
            data_im_in(18)=>mul_im_out(601),
            data_im_in(19)=>mul_im_out(633),
            data_im_in(20)=>mul_im_out(665),
            data_im_in(21)=>mul_im_out(697),
            data_im_in(22)=>mul_im_out(729),
            data_im_in(23)=>mul_im_out(761),
            data_im_in(24)=>mul_im_out(793),
            data_im_in(25)=>mul_im_out(825),
            data_im_in(26)=>mul_im_out(857),
            data_im_in(27)=>mul_im_out(889),
            data_im_in(28)=>mul_im_out(921),
            data_im_in(29)=>mul_im_out(953),
            data_im_in(30)=>mul_im_out(985),
            data_im_in(31)=>mul_im_out(1017),
            data_im_in(32)=>mul_im_out(1049),
            data_im_in(33)=>mul_im_out(1081),
            data_im_in(34)=>mul_im_out(1113),
            data_im_in(35)=>mul_im_out(1145),
            data_im_in(36)=>mul_im_out(1177),
            data_im_in(37)=>mul_im_out(1209),
            data_im_in(38)=>mul_im_out(1241),
            data_im_in(39)=>mul_im_out(1273),
            data_im_in(40)=>mul_im_out(1305),
            data_im_in(41)=>mul_im_out(1337),
            data_im_in(42)=>mul_im_out(1369),
            data_im_in(43)=>mul_im_out(1401),
            data_im_in(44)=>mul_im_out(1433),
            data_im_in(45)=>mul_im_out(1465),
            data_im_in(46)=>mul_im_out(1497),
            data_im_in(47)=>mul_im_out(1529),
            data_im_in(48)=>mul_im_out(1561),
            data_im_in(49)=>mul_im_out(1593),
            data_im_in(50)=>mul_im_out(1625),
            data_im_in(51)=>mul_im_out(1657),
            data_im_in(52)=>mul_im_out(1689),
            data_im_in(53)=>mul_im_out(1721),
            data_im_in(54)=>mul_im_out(1753),
            data_im_in(55)=>mul_im_out(1785),
            data_im_in(56)=>mul_im_out(1817),
            data_im_in(57)=>mul_im_out(1849),
            data_im_in(58)=>mul_im_out(1881),
            data_im_in(59)=>mul_im_out(1913),
            data_im_in(60)=>mul_im_out(1945),
            data_im_in(61)=>mul_im_out(1977),
            data_im_in(62)=>mul_im_out(2009),
            data_im_in(63)=>mul_im_out(2041),
            data_re_out(0)=>data_re_out(25),
            data_re_out(1)=>data_re_out(57),
            data_re_out(2)=>data_re_out(89),
            data_re_out(3)=>data_re_out(121),
            data_re_out(4)=>data_re_out(153),
            data_re_out(5)=>data_re_out(185),
            data_re_out(6)=>data_re_out(217),
            data_re_out(7)=>data_re_out(249),
            data_re_out(8)=>data_re_out(281),
            data_re_out(9)=>data_re_out(313),
            data_re_out(10)=>data_re_out(345),
            data_re_out(11)=>data_re_out(377),
            data_re_out(12)=>data_re_out(409),
            data_re_out(13)=>data_re_out(441),
            data_re_out(14)=>data_re_out(473),
            data_re_out(15)=>data_re_out(505),
            data_re_out(16)=>data_re_out(537),
            data_re_out(17)=>data_re_out(569),
            data_re_out(18)=>data_re_out(601),
            data_re_out(19)=>data_re_out(633),
            data_re_out(20)=>data_re_out(665),
            data_re_out(21)=>data_re_out(697),
            data_re_out(22)=>data_re_out(729),
            data_re_out(23)=>data_re_out(761),
            data_re_out(24)=>data_re_out(793),
            data_re_out(25)=>data_re_out(825),
            data_re_out(26)=>data_re_out(857),
            data_re_out(27)=>data_re_out(889),
            data_re_out(28)=>data_re_out(921),
            data_re_out(29)=>data_re_out(953),
            data_re_out(30)=>data_re_out(985),
            data_re_out(31)=>data_re_out(1017),
            data_re_out(32)=>data_re_out(1049),
            data_re_out(33)=>data_re_out(1081),
            data_re_out(34)=>data_re_out(1113),
            data_re_out(35)=>data_re_out(1145),
            data_re_out(36)=>data_re_out(1177),
            data_re_out(37)=>data_re_out(1209),
            data_re_out(38)=>data_re_out(1241),
            data_re_out(39)=>data_re_out(1273),
            data_re_out(40)=>data_re_out(1305),
            data_re_out(41)=>data_re_out(1337),
            data_re_out(42)=>data_re_out(1369),
            data_re_out(43)=>data_re_out(1401),
            data_re_out(44)=>data_re_out(1433),
            data_re_out(45)=>data_re_out(1465),
            data_re_out(46)=>data_re_out(1497),
            data_re_out(47)=>data_re_out(1529),
            data_re_out(48)=>data_re_out(1561),
            data_re_out(49)=>data_re_out(1593),
            data_re_out(50)=>data_re_out(1625),
            data_re_out(51)=>data_re_out(1657),
            data_re_out(52)=>data_re_out(1689),
            data_re_out(53)=>data_re_out(1721),
            data_re_out(54)=>data_re_out(1753),
            data_re_out(55)=>data_re_out(1785),
            data_re_out(56)=>data_re_out(1817),
            data_re_out(57)=>data_re_out(1849),
            data_re_out(58)=>data_re_out(1881),
            data_re_out(59)=>data_re_out(1913),
            data_re_out(60)=>data_re_out(1945),
            data_re_out(61)=>data_re_out(1977),
            data_re_out(62)=>data_re_out(2009),
            data_re_out(63)=>data_re_out(2041),
            data_im_out(0)=>data_im_out(25),
            data_im_out(1)=>data_im_out(57),
            data_im_out(2)=>data_im_out(89),
            data_im_out(3)=>data_im_out(121),
            data_im_out(4)=>data_im_out(153),
            data_im_out(5)=>data_im_out(185),
            data_im_out(6)=>data_im_out(217),
            data_im_out(7)=>data_im_out(249),
            data_im_out(8)=>data_im_out(281),
            data_im_out(9)=>data_im_out(313),
            data_im_out(10)=>data_im_out(345),
            data_im_out(11)=>data_im_out(377),
            data_im_out(12)=>data_im_out(409),
            data_im_out(13)=>data_im_out(441),
            data_im_out(14)=>data_im_out(473),
            data_im_out(15)=>data_im_out(505),
            data_im_out(16)=>data_im_out(537),
            data_im_out(17)=>data_im_out(569),
            data_im_out(18)=>data_im_out(601),
            data_im_out(19)=>data_im_out(633),
            data_im_out(20)=>data_im_out(665),
            data_im_out(21)=>data_im_out(697),
            data_im_out(22)=>data_im_out(729),
            data_im_out(23)=>data_im_out(761),
            data_im_out(24)=>data_im_out(793),
            data_im_out(25)=>data_im_out(825),
            data_im_out(26)=>data_im_out(857),
            data_im_out(27)=>data_im_out(889),
            data_im_out(28)=>data_im_out(921),
            data_im_out(29)=>data_im_out(953),
            data_im_out(30)=>data_im_out(985),
            data_im_out(31)=>data_im_out(1017),
            data_im_out(32)=>data_im_out(1049),
            data_im_out(33)=>data_im_out(1081),
            data_im_out(34)=>data_im_out(1113),
            data_im_out(35)=>data_im_out(1145),
            data_im_out(36)=>data_im_out(1177),
            data_im_out(37)=>data_im_out(1209),
            data_im_out(38)=>data_im_out(1241),
            data_im_out(39)=>data_im_out(1273),
            data_im_out(40)=>data_im_out(1305),
            data_im_out(41)=>data_im_out(1337),
            data_im_out(42)=>data_im_out(1369),
            data_im_out(43)=>data_im_out(1401),
            data_im_out(44)=>data_im_out(1433),
            data_im_out(45)=>data_im_out(1465),
            data_im_out(46)=>data_im_out(1497),
            data_im_out(47)=>data_im_out(1529),
            data_im_out(48)=>data_im_out(1561),
            data_im_out(49)=>data_im_out(1593),
            data_im_out(50)=>data_im_out(1625),
            data_im_out(51)=>data_im_out(1657),
            data_im_out(52)=>data_im_out(1689),
            data_im_out(53)=>data_im_out(1721),
            data_im_out(54)=>data_im_out(1753),
            data_im_out(55)=>data_im_out(1785),
            data_im_out(56)=>data_im_out(1817),
            data_im_out(57)=>data_im_out(1849),
            data_im_out(58)=>data_im_out(1881),
            data_im_out(59)=>data_im_out(1913),
            data_im_out(60)=>data_im_out(1945),
            data_im_out(61)=>data_im_out(1977),
            data_im_out(62)=>data_im_out(2009),
            data_im_out(63)=>data_im_out(2041)
        );           

    URFFT_PT64_26 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(26),
            data_re_in(1)=>mul_re_out(58),
            data_re_in(2)=>mul_re_out(90),
            data_re_in(3)=>mul_re_out(122),
            data_re_in(4)=>mul_re_out(154),
            data_re_in(5)=>mul_re_out(186),
            data_re_in(6)=>mul_re_out(218),
            data_re_in(7)=>mul_re_out(250),
            data_re_in(8)=>mul_re_out(282),
            data_re_in(9)=>mul_re_out(314),
            data_re_in(10)=>mul_re_out(346),
            data_re_in(11)=>mul_re_out(378),
            data_re_in(12)=>mul_re_out(410),
            data_re_in(13)=>mul_re_out(442),
            data_re_in(14)=>mul_re_out(474),
            data_re_in(15)=>mul_re_out(506),
            data_re_in(16)=>mul_re_out(538),
            data_re_in(17)=>mul_re_out(570),
            data_re_in(18)=>mul_re_out(602),
            data_re_in(19)=>mul_re_out(634),
            data_re_in(20)=>mul_re_out(666),
            data_re_in(21)=>mul_re_out(698),
            data_re_in(22)=>mul_re_out(730),
            data_re_in(23)=>mul_re_out(762),
            data_re_in(24)=>mul_re_out(794),
            data_re_in(25)=>mul_re_out(826),
            data_re_in(26)=>mul_re_out(858),
            data_re_in(27)=>mul_re_out(890),
            data_re_in(28)=>mul_re_out(922),
            data_re_in(29)=>mul_re_out(954),
            data_re_in(30)=>mul_re_out(986),
            data_re_in(31)=>mul_re_out(1018),
            data_re_in(32)=>mul_re_out(1050),
            data_re_in(33)=>mul_re_out(1082),
            data_re_in(34)=>mul_re_out(1114),
            data_re_in(35)=>mul_re_out(1146),
            data_re_in(36)=>mul_re_out(1178),
            data_re_in(37)=>mul_re_out(1210),
            data_re_in(38)=>mul_re_out(1242),
            data_re_in(39)=>mul_re_out(1274),
            data_re_in(40)=>mul_re_out(1306),
            data_re_in(41)=>mul_re_out(1338),
            data_re_in(42)=>mul_re_out(1370),
            data_re_in(43)=>mul_re_out(1402),
            data_re_in(44)=>mul_re_out(1434),
            data_re_in(45)=>mul_re_out(1466),
            data_re_in(46)=>mul_re_out(1498),
            data_re_in(47)=>mul_re_out(1530),
            data_re_in(48)=>mul_re_out(1562),
            data_re_in(49)=>mul_re_out(1594),
            data_re_in(50)=>mul_re_out(1626),
            data_re_in(51)=>mul_re_out(1658),
            data_re_in(52)=>mul_re_out(1690),
            data_re_in(53)=>mul_re_out(1722),
            data_re_in(54)=>mul_re_out(1754),
            data_re_in(55)=>mul_re_out(1786),
            data_re_in(56)=>mul_re_out(1818),
            data_re_in(57)=>mul_re_out(1850),
            data_re_in(58)=>mul_re_out(1882),
            data_re_in(59)=>mul_re_out(1914),
            data_re_in(60)=>mul_re_out(1946),
            data_re_in(61)=>mul_re_out(1978),
            data_re_in(62)=>mul_re_out(2010),
            data_re_in(63)=>mul_re_out(2042),
            data_im_in(0)=>mul_im_out(26),
            data_im_in(1)=>mul_im_out(58),
            data_im_in(2)=>mul_im_out(90),
            data_im_in(3)=>mul_im_out(122),
            data_im_in(4)=>mul_im_out(154),
            data_im_in(5)=>mul_im_out(186),
            data_im_in(6)=>mul_im_out(218),
            data_im_in(7)=>mul_im_out(250),
            data_im_in(8)=>mul_im_out(282),
            data_im_in(9)=>mul_im_out(314),
            data_im_in(10)=>mul_im_out(346),
            data_im_in(11)=>mul_im_out(378),
            data_im_in(12)=>mul_im_out(410),
            data_im_in(13)=>mul_im_out(442),
            data_im_in(14)=>mul_im_out(474),
            data_im_in(15)=>mul_im_out(506),
            data_im_in(16)=>mul_im_out(538),
            data_im_in(17)=>mul_im_out(570),
            data_im_in(18)=>mul_im_out(602),
            data_im_in(19)=>mul_im_out(634),
            data_im_in(20)=>mul_im_out(666),
            data_im_in(21)=>mul_im_out(698),
            data_im_in(22)=>mul_im_out(730),
            data_im_in(23)=>mul_im_out(762),
            data_im_in(24)=>mul_im_out(794),
            data_im_in(25)=>mul_im_out(826),
            data_im_in(26)=>mul_im_out(858),
            data_im_in(27)=>mul_im_out(890),
            data_im_in(28)=>mul_im_out(922),
            data_im_in(29)=>mul_im_out(954),
            data_im_in(30)=>mul_im_out(986),
            data_im_in(31)=>mul_im_out(1018),
            data_im_in(32)=>mul_im_out(1050),
            data_im_in(33)=>mul_im_out(1082),
            data_im_in(34)=>mul_im_out(1114),
            data_im_in(35)=>mul_im_out(1146),
            data_im_in(36)=>mul_im_out(1178),
            data_im_in(37)=>mul_im_out(1210),
            data_im_in(38)=>mul_im_out(1242),
            data_im_in(39)=>mul_im_out(1274),
            data_im_in(40)=>mul_im_out(1306),
            data_im_in(41)=>mul_im_out(1338),
            data_im_in(42)=>mul_im_out(1370),
            data_im_in(43)=>mul_im_out(1402),
            data_im_in(44)=>mul_im_out(1434),
            data_im_in(45)=>mul_im_out(1466),
            data_im_in(46)=>mul_im_out(1498),
            data_im_in(47)=>mul_im_out(1530),
            data_im_in(48)=>mul_im_out(1562),
            data_im_in(49)=>mul_im_out(1594),
            data_im_in(50)=>mul_im_out(1626),
            data_im_in(51)=>mul_im_out(1658),
            data_im_in(52)=>mul_im_out(1690),
            data_im_in(53)=>mul_im_out(1722),
            data_im_in(54)=>mul_im_out(1754),
            data_im_in(55)=>mul_im_out(1786),
            data_im_in(56)=>mul_im_out(1818),
            data_im_in(57)=>mul_im_out(1850),
            data_im_in(58)=>mul_im_out(1882),
            data_im_in(59)=>mul_im_out(1914),
            data_im_in(60)=>mul_im_out(1946),
            data_im_in(61)=>mul_im_out(1978),
            data_im_in(62)=>mul_im_out(2010),
            data_im_in(63)=>mul_im_out(2042),
            data_re_out(0)=>data_re_out(26),
            data_re_out(1)=>data_re_out(58),
            data_re_out(2)=>data_re_out(90),
            data_re_out(3)=>data_re_out(122),
            data_re_out(4)=>data_re_out(154),
            data_re_out(5)=>data_re_out(186),
            data_re_out(6)=>data_re_out(218),
            data_re_out(7)=>data_re_out(250),
            data_re_out(8)=>data_re_out(282),
            data_re_out(9)=>data_re_out(314),
            data_re_out(10)=>data_re_out(346),
            data_re_out(11)=>data_re_out(378),
            data_re_out(12)=>data_re_out(410),
            data_re_out(13)=>data_re_out(442),
            data_re_out(14)=>data_re_out(474),
            data_re_out(15)=>data_re_out(506),
            data_re_out(16)=>data_re_out(538),
            data_re_out(17)=>data_re_out(570),
            data_re_out(18)=>data_re_out(602),
            data_re_out(19)=>data_re_out(634),
            data_re_out(20)=>data_re_out(666),
            data_re_out(21)=>data_re_out(698),
            data_re_out(22)=>data_re_out(730),
            data_re_out(23)=>data_re_out(762),
            data_re_out(24)=>data_re_out(794),
            data_re_out(25)=>data_re_out(826),
            data_re_out(26)=>data_re_out(858),
            data_re_out(27)=>data_re_out(890),
            data_re_out(28)=>data_re_out(922),
            data_re_out(29)=>data_re_out(954),
            data_re_out(30)=>data_re_out(986),
            data_re_out(31)=>data_re_out(1018),
            data_re_out(32)=>data_re_out(1050),
            data_re_out(33)=>data_re_out(1082),
            data_re_out(34)=>data_re_out(1114),
            data_re_out(35)=>data_re_out(1146),
            data_re_out(36)=>data_re_out(1178),
            data_re_out(37)=>data_re_out(1210),
            data_re_out(38)=>data_re_out(1242),
            data_re_out(39)=>data_re_out(1274),
            data_re_out(40)=>data_re_out(1306),
            data_re_out(41)=>data_re_out(1338),
            data_re_out(42)=>data_re_out(1370),
            data_re_out(43)=>data_re_out(1402),
            data_re_out(44)=>data_re_out(1434),
            data_re_out(45)=>data_re_out(1466),
            data_re_out(46)=>data_re_out(1498),
            data_re_out(47)=>data_re_out(1530),
            data_re_out(48)=>data_re_out(1562),
            data_re_out(49)=>data_re_out(1594),
            data_re_out(50)=>data_re_out(1626),
            data_re_out(51)=>data_re_out(1658),
            data_re_out(52)=>data_re_out(1690),
            data_re_out(53)=>data_re_out(1722),
            data_re_out(54)=>data_re_out(1754),
            data_re_out(55)=>data_re_out(1786),
            data_re_out(56)=>data_re_out(1818),
            data_re_out(57)=>data_re_out(1850),
            data_re_out(58)=>data_re_out(1882),
            data_re_out(59)=>data_re_out(1914),
            data_re_out(60)=>data_re_out(1946),
            data_re_out(61)=>data_re_out(1978),
            data_re_out(62)=>data_re_out(2010),
            data_re_out(63)=>data_re_out(2042),
            data_im_out(0)=>data_im_out(26),
            data_im_out(1)=>data_im_out(58),
            data_im_out(2)=>data_im_out(90),
            data_im_out(3)=>data_im_out(122),
            data_im_out(4)=>data_im_out(154),
            data_im_out(5)=>data_im_out(186),
            data_im_out(6)=>data_im_out(218),
            data_im_out(7)=>data_im_out(250),
            data_im_out(8)=>data_im_out(282),
            data_im_out(9)=>data_im_out(314),
            data_im_out(10)=>data_im_out(346),
            data_im_out(11)=>data_im_out(378),
            data_im_out(12)=>data_im_out(410),
            data_im_out(13)=>data_im_out(442),
            data_im_out(14)=>data_im_out(474),
            data_im_out(15)=>data_im_out(506),
            data_im_out(16)=>data_im_out(538),
            data_im_out(17)=>data_im_out(570),
            data_im_out(18)=>data_im_out(602),
            data_im_out(19)=>data_im_out(634),
            data_im_out(20)=>data_im_out(666),
            data_im_out(21)=>data_im_out(698),
            data_im_out(22)=>data_im_out(730),
            data_im_out(23)=>data_im_out(762),
            data_im_out(24)=>data_im_out(794),
            data_im_out(25)=>data_im_out(826),
            data_im_out(26)=>data_im_out(858),
            data_im_out(27)=>data_im_out(890),
            data_im_out(28)=>data_im_out(922),
            data_im_out(29)=>data_im_out(954),
            data_im_out(30)=>data_im_out(986),
            data_im_out(31)=>data_im_out(1018),
            data_im_out(32)=>data_im_out(1050),
            data_im_out(33)=>data_im_out(1082),
            data_im_out(34)=>data_im_out(1114),
            data_im_out(35)=>data_im_out(1146),
            data_im_out(36)=>data_im_out(1178),
            data_im_out(37)=>data_im_out(1210),
            data_im_out(38)=>data_im_out(1242),
            data_im_out(39)=>data_im_out(1274),
            data_im_out(40)=>data_im_out(1306),
            data_im_out(41)=>data_im_out(1338),
            data_im_out(42)=>data_im_out(1370),
            data_im_out(43)=>data_im_out(1402),
            data_im_out(44)=>data_im_out(1434),
            data_im_out(45)=>data_im_out(1466),
            data_im_out(46)=>data_im_out(1498),
            data_im_out(47)=>data_im_out(1530),
            data_im_out(48)=>data_im_out(1562),
            data_im_out(49)=>data_im_out(1594),
            data_im_out(50)=>data_im_out(1626),
            data_im_out(51)=>data_im_out(1658),
            data_im_out(52)=>data_im_out(1690),
            data_im_out(53)=>data_im_out(1722),
            data_im_out(54)=>data_im_out(1754),
            data_im_out(55)=>data_im_out(1786),
            data_im_out(56)=>data_im_out(1818),
            data_im_out(57)=>data_im_out(1850),
            data_im_out(58)=>data_im_out(1882),
            data_im_out(59)=>data_im_out(1914),
            data_im_out(60)=>data_im_out(1946),
            data_im_out(61)=>data_im_out(1978),
            data_im_out(62)=>data_im_out(2010),
            data_im_out(63)=>data_im_out(2042)
        );           

    URFFT_PT64_27 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(27),
            data_re_in(1)=>mul_re_out(59),
            data_re_in(2)=>mul_re_out(91),
            data_re_in(3)=>mul_re_out(123),
            data_re_in(4)=>mul_re_out(155),
            data_re_in(5)=>mul_re_out(187),
            data_re_in(6)=>mul_re_out(219),
            data_re_in(7)=>mul_re_out(251),
            data_re_in(8)=>mul_re_out(283),
            data_re_in(9)=>mul_re_out(315),
            data_re_in(10)=>mul_re_out(347),
            data_re_in(11)=>mul_re_out(379),
            data_re_in(12)=>mul_re_out(411),
            data_re_in(13)=>mul_re_out(443),
            data_re_in(14)=>mul_re_out(475),
            data_re_in(15)=>mul_re_out(507),
            data_re_in(16)=>mul_re_out(539),
            data_re_in(17)=>mul_re_out(571),
            data_re_in(18)=>mul_re_out(603),
            data_re_in(19)=>mul_re_out(635),
            data_re_in(20)=>mul_re_out(667),
            data_re_in(21)=>mul_re_out(699),
            data_re_in(22)=>mul_re_out(731),
            data_re_in(23)=>mul_re_out(763),
            data_re_in(24)=>mul_re_out(795),
            data_re_in(25)=>mul_re_out(827),
            data_re_in(26)=>mul_re_out(859),
            data_re_in(27)=>mul_re_out(891),
            data_re_in(28)=>mul_re_out(923),
            data_re_in(29)=>mul_re_out(955),
            data_re_in(30)=>mul_re_out(987),
            data_re_in(31)=>mul_re_out(1019),
            data_re_in(32)=>mul_re_out(1051),
            data_re_in(33)=>mul_re_out(1083),
            data_re_in(34)=>mul_re_out(1115),
            data_re_in(35)=>mul_re_out(1147),
            data_re_in(36)=>mul_re_out(1179),
            data_re_in(37)=>mul_re_out(1211),
            data_re_in(38)=>mul_re_out(1243),
            data_re_in(39)=>mul_re_out(1275),
            data_re_in(40)=>mul_re_out(1307),
            data_re_in(41)=>mul_re_out(1339),
            data_re_in(42)=>mul_re_out(1371),
            data_re_in(43)=>mul_re_out(1403),
            data_re_in(44)=>mul_re_out(1435),
            data_re_in(45)=>mul_re_out(1467),
            data_re_in(46)=>mul_re_out(1499),
            data_re_in(47)=>mul_re_out(1531),
            data_re_in(48)=>mul_re_out(1563),
            data_re_in(49)=>mul_re_out(1595),
            data_re_in(50)=>mul_re_out(1627),
            data_re_in(51)=>mul_re_out(1659),
            data_re_in(52)=>mul_re_out(1691),
            data_re_in(53)=>mul_re_out(1723),
            data_re_in(54)=>mul_re_out(1755),
            data_re_in(55)=>mul_re_out(1787),
            data_re_in(56)=>mul_re_out(1819),
            data_re_in(57)=>mul_re_out(1851),
            data_re_in(58)=>mul_re_out(1883),
            data_re_in(59)=>mul_re_out(1915),
            data_re_in(60)=>mul_re_out(1947),
            data_re_in(61)=>mul_re_out(1979),
            data_re_in(62)=>mul_re_out(2011),
            data_re_in(63)=>mul_re_out(2043),
            data_im_in(0)=>mul_im_out(27),
            data_im_in(1)=>mul_im_out(59),
            data_im_in(2)=>mul_im_out(91),
            data_im_in(3)=>mul_im_out(123),
            data_im_in(4)=>mul_im_out(155),
            data_im_in(5)=>mul_im_out(187),
            data_im_in(6)=>mul_im_out(219),
            data_im_in(7)=>mul_im_out(251),
            data_im_in(8)=>mul_im_out(283),
            data_im_in(9)=>mul_im_out(315),
            data_im_in(10)=>mul_im_out(347),
            data_im_in(11)=>mul_im_out(379),
            data_im_in(12)=>mul_im_out(411),
            data_im_in(13)=>mul_im_out(443),
            data_im_in(14)=>mul_im_out(475),
            data_im_in(15)=>mul_im_out(507),
            data_im_in(16)=>mul_im_out(539),
            data_im_in(17)=>mul_im_out(571),
            data_im_in(18)=>mul_im_out(603),
            data_im_in(19)=>mul_im_out(635),
            data_im_in(20)=>mul_im_out(667),
            data_im_in(21)=>mul_im_out(699),
            data_im_in(22)=>mul_im_out(731),
            data_im_in(23)=>mul_im_out(763),
            data_im_in(24)=>mul_im_out(795),
            data_im_in(25)=>mul_im_out(827),
            data_im_in(26)=>mul_im_out(859),
            data_im_in(27)=>mul_im_out(891),
            data_im_in(28)=>mul_im_out(923),
            data_im_in(29)=>mul_im_out(955),
            data_im_in(30)=>mul_im_out(987),
            data_im_in(31)=>mul_im_out(1019),
            data_im_in(32)=>mul_im_out(1051),
            data_im_in(33)=>mul_im_out(1083),
            data_im_in(34)=>mul_im_out(1115),
            data_im_in(35)=>mul_im_out(1147),
            data_im_in(36)=>mul_im_out(1179),
            data_im_in(37)=>mul_im_out(1211),
            data_im_in(38)=>mul_im_out(1243),
            data_im_in(39)=>mul_im_out(1275),
            data_im_in(40)=>mul_im_out(1307),
            data_im_in(41)=>mul_im_out(1339),
            data_im_in(42)=>mul_im_out(1371),
            data_im_in(43)=>mul_im_out(1403),
            data_im_in(44)=>mul_im_out(1435),
            data_im_in(45)=>mul_im_out(1467),
            data_im_in(46)=>mul_im_out(1499),
            data_im_in(47)=>mul_im_out(1531),
            data_im_in(48)=>mul_im_out(1563),
            data_im_in(49)=>mul_im_out(1595),
            data_im_in(50)=>mul_im_out(1627),
            data_im_in(51)=>mul_im_out(1659),
            data_im_in(52)=>mul_im_out(1691),
            data_im_in(53)=>mul_im_out(1723),
            data_im_in(54)=>mul_im_out(1755),
            data_im_in(55)=>mul_im_out(1787),
            data_im_in(56)=>mul_im_out(1819),
            data_im_in(57)=>mul_im_out(1851),
            data_im_in(58)=>mul_im_out(1883),
            data_im_in(59)=>mul_im_out(1915),
            data_im_in(60)=>mul_im_out(1947),
            data_im_in(61)=>mul_im_out(1979),
            data_im_in(62)=>mul_im_out(2011),
            data_im_in(63)=>mul_im_out(2043),
            data_re_out(0)=>data_re_out(27),
            data_re_out(1)=>data_re_out(59),
            data_re_out(2)=>data_re_out(91),
            data_re_out(3)=>data_re_out(123),
            data_re_out(4)=>data_re_out(155),
            data_re_out(5)=>data_re_out(187),
            data_re_out(6)=>data_re_out(219),
            data_re_out(7)=>data_re_out(251),
            data_re_out(8)=>data_re_out(283),
            data_re_out(9)=>data_re_out(315),
            data_re_out(10)=>data_re_out(347),
            data_re_out(11)=>data_re_out(379),
            data_re_out(12)=>data_re_out(411),
            data_re_out(13)=>data_re_out(443),
            data_re_out(14)=>data_re_out(475),
            data_re_out(15)=>data_re_out(507),
            data_re_out(16)=>data_re_out(539),
            data_re_out(17)=>data_re_out(571),
            data_re_out(18)=>data_re_out(603),
            data_re_out(19)=>data_re_out(635),
            data_re_out(20)=>data_re_out(667),
            data_re_out(21)=>data_re_out(699),
            data_re_out(22)=>data_re_out(731),
            data_re_out(23)=>data_re_out(763),
            data_re_out(24)=>data_re_out(795),
            data_re_out(25)=>data_re_out(827),
            data_re_out(26)=>data_re_out(859),
            data_re_out(27)=>data_re_out(891),
            data_re_out(28)=>data_re_out(923),
            data_re_out(29)=>data_re_out(955),
            data_re_out(30)=>data_re_out(987),
            data_re_out(31)=>data_re_out(1019),
            data_re_out(32)=>data_re_out(1051),
            data_re_out(33)=>data_re_out(1083),
            data_re_out(34)=>data_re_out(1115),
            data_re_out(35)=>data_re_out(1147),
            data_re_out(36)=>data_re_out(1179),
            data_re_out(37)=>data_re_out(1211),
            data_re_out(38)=>data_re_out(1243),
            data_re_out(39)=>data_re_out(1275),
            data_re_out(40)=>data_re_out(1307),
            data_re_out(41)=>data_re_out(1339),
            data_re_out(42)=>data_re_out(1371),
            data_re_out(43)=>data_re_out(1403),
            data_re_out(44)=>data_re_out(1435),
            data_re_out(45)=>data_re_out(1467),
            data_re_out(46)=>data_re_out(1499),
            data_re_out(47)=>data_re_out(1531),
            data_re_out(48)=>data_re_out(1563),
            data_re_out(49)=>data_re_out(1595),
            data_re_out(50)=>data_re_out(1627),
            data_re_out(51)=>data_re_out(1659),
            data_re_out(52)=>data_re_out(1691),
            data_re_out(53)=>data_re_out(1723),
            data_re_out(54)=>data_re_out(1755),
            data_re_out(55)=>data_re_out(1787),
            data_re_out(56)=>data_re_out(1819),
            data_re_out(57)=>data_re_out(1851),
            data_re_out(58)=>data_re_out(1883),
            data_re_out(59)=>data_re_out(1915),
            data_re_out(60)=>data_re_out(1947),
            data_re_out(61)=>data_re_out(1979),
            data_re_out(62)=>data_re_out(2011),
            data_re_out(63)=>data_re_out(2043),
            data_im_out(0)=>data_im_out(27),
            data_im_out(1)=>data_im_out(59),
            data_im_out(2)=>data_im_out(91),
            data_im_out(3)=>data_im_out(123),
            data_im_out(4)=>data_im_out(155),
            data_im_out(5)=>data_im_out(187),
            data_im_out(6)=>data_im_out(219),
            data_im_out(7)=>data_im_out(251),
            data_im_out(8)=>data_im_out(283),
            data_im_out(9)=>data_im_out(315),
            data_im_out(10)=>data_im_out(347),
            data_im_out(11)=>data_im_out(379),
            data_im_out(12)=>data_im_out(411),
            data_im_out(13)=>data_im_out(443),
            data_im_out(14)=>data_im_out(475),
            data_im_out(15)=>data_im_out(507),
            data_im_out(16)=>data_im_out(539),
            data_im_out(17)=>data_im_out(571),
            data_im_out(18)=>data_im_out(603),
            data_im_out(19)=>data_im_out(635),
            data_im_out(20)=>data_im_out(667),
            data_im_out(21)=>data_im_out(699),
            data_im_out(22)=>data_im_out(731),
            data_im_out(23)=>data_im_out(763),
            data_im_out(24)=>data_im_out(795),
            data_im_out(25)=>data_im_out(827),
            data_im_out(26)=>data_im_out(859),
            data_im_out(27)=>data_im_out(891),
            data_im_out(28)=>data_im_out(923),
            data_im_out(29)=>data_im_out(955),
            data_im_out(30)=>data_im_out(987),
            data_im_out(31)=>data_im_out(1019),
            data_im_out(32)=>data_im_out(1051),
            data_im_out(33)=>data_im_out(1083),
            data_im_out(34)=>data_im_out(1115),
            data_im_out(35)=>data_im_out(1147),
            data_im_out(36)=>data_im_out(1179),
            data_im_out(37)=>data_im_out(1211),
            data_im_out(38)=>data_im_out(1243),
            data_im_out(39)=>data_im_out(1275),
            data_im_out(40)=>data_im_out(1307),
            data_im_out(41)=>data_im_out(1339),
            data_im_out(42)=>data_im_out(1371),
            data_im_out(43)=>data_im_out(1403),
            data_im_out(44)=>data_im_out(1435),
            data_im_out(45)=>data_im_out(1467),
            data_im_out(46)=>data_im_out(1499),
            data_im_out(47)=>data_im_out(1531),
            data_im_out(48)=>data_im_out(1563),
            data_im_out(49)=>data_im_out(1595),
            data_im_out(50)=>data_im_out(1627),
            data_im_out(51)=>data_im_out(1659),
            data_im_out(52)=>data_im_out(1691),
            data_im_out(53)=>data_im_out(1723),
            data_im_out(54)=>data_im_out(1755),
            data_im_out(55)=>data_im_out(1787),
            data_im_out(56)=>data_im_out(1819),
            data_im_out(57)=>data_im_out(1851),
            data_im_out(58)=>data_im_out(1883),
            data_im_out(59)=>data_im_out(1915),
            data_im_out(60)=>data_im_out(1947),
            data_im_out(61)=>data_im_out(1979),
            data_im_out(62)=>data_im_out(2011),
            data_im_out(63)=>data_im_out(2043)
        );           

    URFFT_PT64_28 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(28),
            data_re_in(1)=>mul_re_out(60),
            data_re_in(2)=>mul_re_out(92),
            data_re_in(3)=>mul_re_out(124),
            data_re_in(4)=>mul_re_out(156),
            data_re_in(5)=>mul_re_out(188),
            data_re_in(6)=>mul_re_out(220),
            data_re_in(7)=>mul_re_out(252),
            data_re_in(8)=>mul_re_out(284),
            data_re_in(9)=>mul_re_out(316),
            data_re_in(10)=>mul_re_out(348),
            data_re_in(11)=>mul_re_out(380),
            data_re_in(12)=>mul_re_out(412),
            data_re_in(13)=>mul_re_out(444),
            data_re_in(14)=>mul_re_out(476),
            data_re_in(15)=>mul_re_out(508),
            data_re_in(16)=>mul_re_out(540),
            data_re_in(17)=>mul_re_out(572),
            data_re_in(18)=>mul_re_out(604),
            data_re_in(19)=>mul_re_out(636),
            data_re_in(20)=>mul_re_out(668),
            data_re_in(21)=>mul_re_out(700),
            data_re_in(22)=>mul_re_out(732),
            data_re_in(23)=>mul_re_out(764),
            data_re_in(24)=>mul_re_out(796),
            data_re_in(25)=>mul_re_out(828),
            data_re_in(26)=>mul_re_out(860),
            data_re_in(27)=>mul_re_out(892),
            data_re_in(28)=>mul_re_out(924),
            data_re_in(29)=>mul_re_out(956),
            data_re_in(30)=>mul_re_out(988),
            data_re_in(31)=>mul_re_out(1020),
            data_re_in(32)=>mul_re_out(1052),
            data_re_in(33)=>mul_re_out(1084),
            data_re_in(34)=>mul_re_out(1116),
            data_re_in(35)=>mul_re_out(1148),
            data_re_in(36)=>mul_re_out(1180),
            data_re_in(37)=>mul_re_out(1212),
            data_re_in(38)=>mul_re_out(1244),
            data_re_in(39)=>mul_re_out(1276),
            data_re_in(40)=>mul_re_out(1308),
            data_re_in(41)=>mul_re_out(1340),
            data_re_in(42)=>mul_re_out(1372),
            data_re_in(43)=>mul_re_out(1404),
            data_re_in(44)=>mul_re_out(1436),
            data_re_in(45)=>mul_re_out(1468),
            data_re_in(46)=>mul_re_out(1500),
            data_re_in(47)=>mul_re_out(1532),
            data_re_in(48)=>mul_re_out(1564),
            data_re_in(49)=>mul_re_out(1596),
            data_re_in(50)=>mul_re_out(1628),
            data_re_in(51)=>mul_re_out(1660),
            data_re_in(52)=>mul_re_out(1692),
            data_re_in(53)=>mul_re_out(1724),
            data_re_in(54)=>mul_re_out(1756),
            data_re_in(55)=>mul_re_out(1788),
            data_re_in(56)=>mul_re_out(1820),
            data_re_in(57)=>mul_re_out(1852),
            data_re_in(58)=>mul_re_out(1884),
            data_re_in(59)=>mul_re_out(1916),
            data_re_in(60)=>mul_re_out(1948),
            data_re_in(61)=>mul_re_out(1980),
            data_re_in(62)=>mul_re_out(2012),
            data_re_in(63)=>mul_re_out(2044),
            data_im_in(0)=>mul_im_out(28),
            data_im_in(1)=>mul_im_out(60),
            data_im_in(2)=>mul_im_out(92),
            data_im_in(3)=>mul_im_out(124),
            data_im_in(4)=>mul_im_out(156),
            data_im_in(5)=>mul_im_out(188),
            data_im_in(6)=>mul_im_out(220),
            data_im_in(7)=>mul_im_out(252),
            data_im_in(8)=>mul_im_out(284),
            data_im_in(9)=>mul_im_out(316),
            data_im_in(10)=>mul_im_out(348),
            data_im_in(11)=>mul_im_out(380),
            data_im_in(12)=>mul_im_out(412),
            data_im_in(13)=>mul_im_out(444),
            data_im_in(14)=>mul_im_out(476),
            data_im_in(15)=>mul_im_out(508),
            data_im_in(16)=>mul_im_out(540),
            data_im_in(17)=>mul_im_out(572),
            data_im_in(18)=>mul_im_out(604),
            data_im_in(19)=>mul_im_out(636),
            data_im_in(20)=>mul_im_out(668),
            data_im_in(21)=>mul_im_out(700),
            data_im_in(22)=>mul_im_out(732),
            data_im_in(23)=>mul_im_out(764),
            data_im_in(24)=>mul_im_out(796),
            data_im_in(25)=>mul_im_out(828),
            data_im_in(26)=>mul_im_out(860),
            data_im_in(27)=>mul_im_out(892),
            data_im_in(28)=>mul_im_out(924),
            data_im_in(29)=>mul_im_out(956),
            data_im_in(30)=>mul_im_out(988),
            data_im_in(31)=>mul_im_out(1020),
            data_im_in(32)=>mul_im_out(1052),
            data_im_in(33)=>mul_im_out(1084),
            data_im_in(34)=>mul_im_out(1116),
            data_im_in(35)=>mul_im_out(1148),
            data_im_in(36)=>mul_im_out(1180),
            data_im_in(37)=>mul_im_out(1212),
            data_im_in(38)=>mul_im_out(1244),
            data_im_in(39)=>mul_im_out(1276),
            data_im_in(40)=>mul_im_out(1308),
            data_im_in(41)=>mul_im_out(1340),
            data_im_in(42)=>mul_im_out(1372),
            data_im_in(43)=>mul_im_out(1404),
            data_im_in(44)=>mul_im_out(1436),
            data_im_in(45)=>mul_im_out(1468),
            data_im_in(46)=>mul_im_out(1500),
            data_im_in(47)=>mul_im_out(1532),
            data_im_in(48)=>mul_im_out(1564),
            data_im_in(49)=>mul_im_out(1596),
            data_im_in(50)=>mul_im_out(1628),
            data_im_in(51)=>mul_im_out(1660),
            data_im_in(52)=>mul_im_out(1692),
            data_im_in(53)=>mul_im_out(1724),
            data_im_in(54)=>mul_im_out(1756),
            data_im_in(55)=>mul_im_out(1788),
            data_im_in(56)=>mul_im_out(1820),
            data_im_in(57)=>mul_im_out(1852),
            data_im_in(58)=>mul_im_out(1884),
            data_im_in(59)=>mul_im_out(1916),
            data_im_in(60)=>mul_im_out(1948),
            data_im_in(61)=>mul_im_out(1980),
            data_im_in(62)=>mul_im_out(2012),
            data_im_in(63)=>mul_im_out(2044),
            data_re_out(0)=>data_re_out(28),
            data_re_out(1)=>data_re_out(60),
            data_re_out(2)=>data_re_out(92),
            data_re_out(3)=>data_re_out(124),
            data_re_out(4)=>data_re_out(156),
            data_re_out(5)=>data_re_out(188),
            data_re_out(6)=>data_re_out(220),
            data_re_out(7)=>data_re_out(252),
            data_re_out(8)=>data_re_out(284),
            data_re_out(9)=>data_re_out(316),
            data_re_out(10)=>data_re_out(348),
            data_re_out(11)=>data_re_out(380),
            data_re_out(12)=>data_re_out(412),
            data_re_out(13)=>data_re_out(444),
            data_re_out(14)=>data_re_out(476),
            data_re_out(15)=>data_re_out(508),
            data_re_out(16)=>data_re_out(540),
            data_re_out(17)=>data_re_out(572),
            data_re_out(18)=>data_re_out(604),
            data_re_out(19)=>data_re_out(636),
            data_re_out(20)=>data_re_out(668),
            data_re_out(21)=>data_re_out(700),
            data_re_out(22)=>data_re_out(732),
            data_re_out(23)=>data_re_out(764),
            data_re_out(24)=>data_re_out(796),
            data_re_out(25)=>data_re_out(828),
            data_re_out(26)=>data_re_out(860),
            data_re_out(27)=>data_re_out(892),
            data_re_out(28)=>data_re_out(924),
            data_re_out(29)=>data_re_out(956),
            data_re_out(30)=>data_re_out(988),
            data_re_out(31)=>data_re_out(1020),
            data_re_out(32)=>data_re_out(1052),
            data_re_out(33)=>data_re_out(1084),
            data_re_out(34)=>data_re_out(1116),
            data_re_out(35)=>data_re_out(1148),
            data_re_out(36)=>data_re_out(1180),
            data_re_out(37)=>data_re_out(1212),
            data_re_out(38)=>data_re_out(1244),
            data_re_out(39)=>data_re_out(1276),
            data_re_out(40)=>data_re_out(1308),
            data_re_out(41)=>data_re_out(1340),
            data_re_out(42)=>data_re_out(1372),
            data_re_out(43)=>data_re_out(1404),
            data_re_out(44)=>data_re_out(1436),
            data_re_out(45)=>data_re_out(1468),
            data_re_out(46)=>data_re_out(1500),
            data_re_out(47)=>data_re_out(1532),
            data_re_out(48)=>data_re_out(1564),
            data_re_out(49)=>data_re_out(1596),
            data_re_out(50)=>data_re_out(1628),
            data_re_out(51)=>data_re_out(1660),
            data_re_out(52)=>data_re_out(1692),
            data_re_out(53)=>data_re_out(1724),
            data_re_out(54)=>data_re_out(1756),
            data_re_out(55)=>data_re_out(1788),
            data_re_out(56)=>data_re_out(1820),
            data_re_out(57)=>data_re_out(1852),
            data_re_out(58)=>data_re_out(1884),
            data_re_out(59)=>data_re_out(1916),
            data_re_out(60)=>data_re_out(1948),
            data_re_out(61)=>data_re_out(1980),
            data_re_out(62)=>data_re_out(2012),
            data_re_out(63)=>data_re_out(2044),
            data_im_out(0)=>data_im_out(28),
            data_im_out(1)=>data_im_out(60),
            data_im_out(2)=>data_im_out(92),
            data_im_out(3)=>data_im_out(124),
            data_im_out(4)=>data_im_out(156),
            data_im_out(5)=>data_im_out(188),
            data_im_out(6)=>data_im_out(220),
            data_im_out(7)=>data_im_out(252),
            data_im_out(8)=>data_im_out(284),
            data_im_out(9)=>data_im_out(316),
            data_im_out(10)=>data_im_out(348),
            data_im_out(11)=>data_im_out(380),
            data_im_out(12)=>data_im_out(412),
            data_im_out(13)=>data_im_out(444),
            data_im_out(14)=>data_im_out(476),
            data_im_out(15)=>data_im_out(508),
            data_im_out(16)=>data_im_out(540),
            data_im_out(17)=>data_im_out(572),
            data_im_out(18)=>data_im_out(604),
            data_im_out(19)=>data_im_out(636),
            data_im_out(20)=>data_im_out(668),
            data_im_out(21)=>data_im_out(700),
            data_im_out(22)=>data_im_out(732),
            data_im_out(23)=>data_im_out(764),
            data_im_out(24)=>data_im_out(796),
            data_im_out(25)=>data_im_out(828),
            data_im_out(26)=>data_im_out(860),
            data_im_out(27)=>data_im_out(892),
            data_im_out(28)=>data_im_out(924),
            data_im_out(29)=>data_im_out(956),
            data_im_out(30)=>data_im_out(988),
            data_im_out(31)=>data_im_out(1020),
            data_im_out(32)=>data_im_out(1052),
            data_im_out(33)=>data_im_out(1084),
            data_im_out(34)=>data_im_out(1116),
            data_im_out(35)=>data_im_out(1148),
            data_im_out(36)=>data_im_out(1180),
            data_im_out(37)=>data_im_out(1212),
            data_im_out(38)=>data_im_out(1244),
            data_im_out(39)=>data_im_out(1276),
            data_im_out(40)=>data_im_out(1308),
            data_im_out(41)=>data_im_out(1340),
            data_im_out(42)=>data_im_out(1372),
            data_im_out(43)=>data_im_out(1404),
            data_im_out(44)=>data_im_out(1436),
            data_im_out(45)=>data_im_out(1468),
            data_im_out(46)=>data_im_out(1500),
            data_im_out(47)=>data_im_out(1532),
            data_im_out(48)=>data_im_out(1564),
            data_im_out(49)=>data_im_out(1596),
            data_im_out(50)=>data_im_out(1628),
            data_im_out(51)=>data_im_out(1660),
            data_im_out(52)=>data_im_out(1692),
            data_im_out(53)=>data_im_out(1724),
            data_im_out(54)=>data_im_out(1756),
            data_im_out(55)=>data_im_out(1788),
            data_im_out(56)=>data_im_out(1820),
            data_im_out(57)=>data_im_out(1852),
            data_im_out(58)=>data_im_out(1884),
            data_im_out(59)=>data_im_out(1916),
            data_im_out(60)=>data_im_out(1948),
            data_im_out(61)=>data_im_out(1980),
            data_im_out(62)=>data_im_out(2012),
            data_im_out(63)=>data_im_out(2044)
        );           

    URFFT_PT64_29 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(29),
            data_re_in(1)=>mul_re_out(61),
            data_re_in(2)=>mul_re_out(93),
            data_re_in(3)=>mul_re_out(125),
            data_re_in(4)=>mul_re_out(157),
            data_re_in(5)=>mul_re_out(189),
            data_re_in(6)=>mul_re_out(221),
            data_re_in(7)=>mul_re_out(253),
            data_re_in(8)=>mul_re_out(285),
            data_re_in(9)=>mul_re_out(317),
            data_re_in(10)=>mul_re_out(349),
            data_re_in(11)=>mul_re_out(381),
            data_re_in(12)=>mul_re_out(413),
            data_re_in(13)=>mul_re_out(445),
            data_re_in(14)=>mul_re_out(477),
            data_re_in(15)=>mul_re_out(509),
            data_re_in(16)=>mul_re_out(541),
            data_re_in(17)=>mul_re_out(573),
            data_re_in(18)=>mul_re_out(605),
            data_re_in(19)=>mul_re_out(637),
            data_re_in(20)=>mul_re_out(669),
            data_re_in(21)=>mul_re_out(701),
            data_re_in(22)=>mul_re_out(733),
            data_re_in(23)=>mul_re_out(765),
            data_re_in(24)=>mul_re_out(797),
            data_re_in(25)=>mul_re_out(829),
            data_re_in(26)=>mul_re_out(861),
            data_re_in(27)=>mul_re_out(893),
            data_re_in(28)=>mul_re_out(925),
            data_re_in(29)=>mul_re_out(957),
            data_re_in(30)=>mul_re_out(989),
            data_re_in(31)=>mul_re_out(1021),
            data_re_in(32)=>mul_re_out(1053),
            data_re_in(33)=>mul_re_out(1085),
            data_re_in(34)=>mul_re_out(1117),
            data_re_in(35)=>mul_re_out(1149),
            data_re_in(36)=>mul_re_out(1181),
            data_re_in(37)=>mul_re_out(1213),
            data_re_in(38)=>mul_re_out(1245),
            data_re_in(39)=>mul_re_out(1277),
            data_re_in(40)=>mul_re_out(1309),
            data_re_in(41)=>mul_re_out(1341),
            data_re_in(42)=>mul_re_out(1373),
            data_re_in(43)=>mul_re_out(1405),
            data_re_in(44)=>mul_re_out(1437),
            data_re_in(45)=>mul_re_out(1469),
            data_re_in(46)=>mul_re_out(1501),
            data_re_in(47)=>mul_re_out(1533),
            data_re_in(48)=>mul_re_out(1565),
            data_re_in(49)=>mul_re_out(1597),
            data_re_in(50)=>mul_re_out(1629),
            data_re_in(51)=>mul_re_out(1661),
            data_re_in(52)=>mul_re_out(1693),
            data_re_in(53)=>mul_re_out(1725),
            data_re_in(54)=>mul_re_out(1757),
            data_re_in(55)=>mul_re_out(1789),
            data_re_in(56)=>mul_re_out(1821),
            data_re_in(57)=>mul_re_out(1853),
            data_re_in(58)=>mul_re_out(1885),
            data_re_in(59)=>mul_re_out(1917),
            data_re_in(60)=>mul_re_out(1949),
            data_re_in(61)=>mul_re_out(1981),
            data_re_in(62)=>mul_re_out(2013),
            data_re_in(63)=>mul_re_out(2045),
            data_im_in(0)=>mul_im_out(29),
            data_im_in(1)=>mul_im_out(61),
            data_im_in(2)=>mul_im_out(93),
            data_im_in(3)=>mul_im_out(125),
            data_im_in(4)=>mul_im_out(157),
            data_im_in(5)=>mul_im_out(189),
            data_im_in(6)=>mul_im_out(221),
            data_im_in(7)=>mul_im_out(253),
            data_im_in(8)=>mul_im_out(285),
            data_im_in(9)=>mul_im_out(317),
            data_im_in(10)=>mul_im_out(349),
            data_im_in(11)=>mul_im_out(381),
            data_im_in(12)=>mul_im_out(413),
            data_im_in(13)=>mul_im_out(445),
            data_im_in(14)=>mul_im_out(477),
            data_im_in(15)=>mul_im_out(509),
            data_im_in(16)=>mul_im_out(541),
            data_im_in(17)=>mul_im_out(573),
            data_im_in(18)=>mul_im_out(605),
            data_im_in(19)=>mul_im_out(637),
            data_im_in(20)=>mul_im_out(669),
            data_im_in(21)=>mul_im_out(701),
            data_im_in(22)=>mul_im_out(733),
            data_im_in(23)=>mul_im_out(765),
            data_im_in(24)=>mul_im_out(797),
            data_im_in(25)=>mul_im_out(829),
            data_im_in(26)=>mul_im_out(861),
            data_im_in(27)=>mul_im_out(893),
            data_im_in(28)=>mul_im_out(925),
            data_im_in(29)=>mul_im_out(957),
            data_im_in(30)=>mul_im_out(989),
            data_im_in(31)=>mul_im_out(1021),
            data_im_in(32)=>mul_im_out(1053),
            data_im_in(33)=>mul_im_out(1085),
            data_im_in(34)=>mul_im_out(1117),
            data_im_in(35)=>mul_im_out(1149),
            data_im_in(36)=>mul_im_out(1181),
            data_im_in(37)=>mul_im_out(1213),
            data_im_in(38)=>mul_im_out(1245),
            data_im_in(39)=>mul_im_out(1277),
            data_im_in(40)=>mul_im_out(1309),
            data_im_in(41)=>mul_im_out(1341),
            data_im_in(42)=>mul_im_out(1373),
            data_im_in(43)=>mul_im_out(1405),
            data_im_in(44)=>mul_im_out(1437),
            data_im_in(45)=>mul_im_out(1469),
            data_im_in(46)=>mul_im_out(1501),
            data_im_in(47)=>mul_im_out(1533),
            data_im_in(48)=>mul_im_out(1565),
            data_im_in(49)=>mul_im_out(1597),
            data_im_in(50)=>mul_im_out(1629),
            data_im_in(51)=>mul_im_out(1661),
            data_im_in(52)=>mul_im_out(1693),
            data_im_in(53)=>mul_im_out(1725),
            data_im_in(54)=>mul_im_out(1757),
            data_im_in(55)=>mul_im_out(1789),
            data_im_in(56)=>mul_im_out(1821),
            data_im_in(57)=>mul_im_out(1853),
            data_im_in(58)=>mul_im_out(1885),
            data_im_in(59)=>mul_im_out(1917),
            data_im_in(60)=>mul_im_out(1949),
            data_im_in(61)=>mul_im_out(1981),
            data_im_in(62)=>mul_im_out(2013),
            data_im_in(63)=>mul_im_out(2045),
            data_re_out(0)=>data_re_out(29),
            data_re_out(1)=>data_re_out(61),
            data_re_out(2)=>data_re_out(93),
            data_re_out(3)=>data_re_out(125),
            data_re_out(4)=>data_re_out(157),
            data_re_out(5)=>data_re_out(189),
            data_re_out(6)=>data_re_out(221),
            data_re_out(7)=>data_re_out(253),
            data_re_out(8)=>data_re_out(285),
            data_re_out(9)=>data_re_out(317),
            data_re_out(10)=>data_re_out(349),
            data_re_out(11)=>data_re_out(381),
            data_re_out(12)=>data_re_out(413),
            data_re_out(13)=>data_re_out(445),
            data_re_out(14)=>data_re_out(477),
            data_re_out(15)=>data_re_out(509),
            data_re_out(16)=>data_re_out(541),
            data_re_out(17)=>data_re_out(573),
            data_re_out(18)=>data_re_out(605),
            data_re_out(19)=>data_re_out(637),
            data_re_out(20)=>data_re_out(669),
            data_re_out(21)=>data_re_out(701),
            data_re_out(22)=>data_re_out(733),
            data_re_out(23)=>data_re_out(765),
            data_re_out(24)=>data_re_out(797),
            data_re_out(25)=>data_re_out(829),
            data_re_out(26)=>data_re_out(861),
            data_re_out(27)=>data_re_out(893),
            data_re_out(28)=>data_re_out(925),
            data_re_out(29)=>data_re_out(957),
            data_re_out(30)=>data_re_out(989),
            data_re_out(31)=>data_re_out(1021),
            data_re_out(32)=>data_re_out(1053),
            data_re_out(33)=>data_re_out(1085),
            data_re_out(34)=>data_re_out(1117),
            data_re_out(35)=>data_re_out(1149),
            data_re_out(36)=>data_re_out(1181),
            data_re_out(37)=>data_re_out(1213),
            data_re_out(38)=>data_re_out(1245),
            data_re_out(39)=>data_re_out(1277),
            data_re_out(40)=>data_re_out(1309),
            data_re_out(41)=>data_re_out(1341),
            data_re_out(42)=>data_re_out(1373),
            data_re_out(43)=>data_re_out(1405),
            data_re_out(44)=>data_re_out(1437),
            data_re_out(45)=>data_re_out(1469),
            data_re_out(46)=>data_re_out(1501),
            data_re_out(47)=>data_re_out(1533),
            data_re_out(48)=>data_re_out(1565),
            data_re_out(49)=>data_re_out(1597),
            data_re_out(50)=>data_re_out(1629),
            data_re_out(51)=>data_re_out(1661),
            data_re_out(52)=>data_re_out(1693),
            data_re_out(53)=>data_re_out(1725),
            data_re_out(54)=>data_re_out(1757),
            data_re_out(55)=>data_re_out(1789),
            data_re_out(56)=>data_re_out(1821),
            data_re_out(57)=>data_re_out(1853),
            data_re_out(58)=>data_re_out(1885),
            data_re_out(59)=>data_re_out(1917),
            data_re_out(60)=>data_re_out(1949),
            data_re_out(61)=>data_re_out(1981),
            data_re_out(62)=>data_re_out(2013),
            data_re_out(63)=>data_re_out(2045),
            data_im_out(0)=>data_im_out(29),
            data_im_out(1)=>data_im_out(61),
            data_im_out(2)=>data_im_out(93),
            data_im_out(3)=>data_im_out(125),
            data_im_out(4)=>data_im_out(157),
            data_im_out(5)=>data_im_out(189),
            data_im_out(6)=>data_im_out(221),
            data_im_out(7)=>data_im_out(253),
            data_im_out(8)=>data_im_out(285),
            data_im_out(9)=>data_im_out(317),
            data_im_out(10)=>data_im_out(349),
            data_im_out(11)=>data_im_out(381),
            data_im_out(12)=>data_im_out(413),
            data_im_out(13)=>data_im_out(445),
            data_im_out(14)=>data_im_out(477),
            data_im_out(15)=>data_im_out(509),
            data_im_out(16)=>data_im_out(541),
            data_im_out(17)=>data_im_out(573),
            data_im_out(18)=>data_im_out(605),
            data_im_out(19)=>data_im_out(637),
            data_im_out(20)=>data_im_out(669),
            data_im_out(21)=>data_im_out(701),
            data_im_out(22)=>data_im_out(733),
            data_im_out(23)=>data_im_out(765),
            data_im_out(24)=>data_im_out(797),
            data_im_out(25)=>data_im_out(829),
            data_im_out(26)=>data_im_out(861),
            data_im_out(27)=>data_im_out(893),
            data_im_out(28)=>data_im_out(925),
            data_im_out(29)=>data_im_out(957),
            data_im_out(30)=>data_im_out(989),
            data_im_out(31)=>data_im_out(1021),
            data_im_out(32)=>data_im_out(1053),
            data_im_out(33)=>data_im_out(1085),
            data_im_out(34)=>data_im_out(1117),
            data_im_out(35)=>data_im_out(1149),
            data_im_out(36)=>data_im_out(1181),
            data_im_out(37)=>data_im_out(1213),
            data_im_out(38)=>data_im_out(1245),
            data_im_out(39)=>data_im_out(1277),
            data_im_out(40)=>data_im_out(1309),
            data_im_out(41)=>data_im_out(1341),
            data_im_out(42)=>data_im_out(1373),
            data_im_out(43)=>data_im_out(1405),
            data_im_out(44)=>data_im_out(1437),
            data_im_out(45)=>data_im_out(1469),
            data_im_out(46)=>data_im_out(1501),
            data_im_out(47)=>data_im_out(1533),
            data_im_out(48)=>data_im_out(1565),
            data_im_out(49)=>data_im_out(1597),
            data_im_out(50)=>data_im_out(1629),
            data_im_out(51)=>data_im_out(1661),
            data_im_out(52)=>data_im_out(1693),
            data_im_out(53)=>data_im_out(1725),
            data_im_out(54)=>data_im_out(1757),
            data_im_out(55)=>data_im_out(1789),
            data_im_out(56)=>data_im_out(1821),
            data_im_out(57)=>data_im_out(1853),
            data_im_out(58)=>data_im_out(1885),
            data_im_out(59)=>data_im_out(1917),
            data_im_out(60)=>data_im_out(1949),
            data_im_out(61)=>data_im_out(1981),
            data_im_out(62)=>data_im_out(2013),
            data_im_out(63)=>data_im_out(2045)
        );           

    URFFT_PT64_30 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(30),
            data_re_in(1)=>mul_re_out(62),
            data_re_in(2)=>mul_re_out(94),
            data_re_in(3)=>mul_re_out(126),
            data_re_in(4)=>mul_re_out(158),
            data_re_in(5)=>mul_re_out(190),
            data_re_in(6)=>mul_re_out(222),
            data_re_in(7)=>mul_re_out(254),
            data_re_in(8)=>mul_re_out(286),
            data_re_in(9)=>mul_re_out(318),
            data_re_in(10)=>mul_re_out(350),
            data_re_in(11)=>mul_re_out(382),
            data_re_in(12)=>mul_re_out(414),
            data_re_in(13)=>mul_re_out(446),
            data_re_in(14)=>mul_re_out(478),
            data_re_in(15)=>mul_re_out(510),
            data_re_in(16)=>mul_re_out(542),
            data_re_in(17)=>mul_re_out(574),
            data_re_in(18)=>mul_re_out(606),
            data_re_in(19)=>mul_re_out(638),
            data_re_in(20)=>mul_re_out(670),
            data_re_in(21)=>mul_re_out(702),
            data_re_in(22)=>mul_re_out(734),
            data_re_in(23)=>mul_re_out(766),
            data_re_in(24)=>mul_re_out(798),
            data_re_in(25)=>mul_re_out(830),
            data_re_in(26)=>mul_re_out(862),
            data_re_in(27)=>mul_re_out(894),
            data_re_in(28)=>mul_re_out(926),
            data_re_in(29)=>mul_re_out(958),
            data_re_in(30)=>mul_re_out(990),
            data_re_in(31)=>mul_re_out(1022),
            data_re_in(32)=>mul_re_out(1054),
            data_re_in(33)=>mul_re_out(1086),
            data_re_in(34)=>mul_re_out(1118),
            data_re_in(35)=>mul_re_out(1150),
            data_re_in(36)=>mul_re_out(1182),
            data_re_in(37)=>mul_re_out(1214),
            data_re_in(38)=>mul_re_out(1246),
            data_re_in(39)=>mul_re_out(1278),
            data_re_in(40)=>mul_re_out(1310),
            data_re_in(41)=>mul_re_out(1342),
            data_re_in(42)=>mul_re_out(1374),
            data_re_in(43)=>mul_re_out(1406),
            data_re_in(44)=>mul_re_out(1438),
            data_re_in(45)=>mul_re_out(1470),
            data_re_in(46)=>mul_re_out(1502),
            data_re_in(47)=>mul_re_out(1534),
            data_re_in(48)=>mul_re_out(1566),
            data_re_in(49)=>mul_re_out(1598),
            data_re_in(50)=>mul_re_out(1630),
            data_re_in(51)=>mul_re_out(1662),
            data_re_in(52)=>mul_re_out(1694),
            data_re_in(53)=>mul_re_out(1726),
            data_re_in(54)=>mul_re_out(1758),
            data_re_in(55)=>mul_re_out(1790),
            data_re_in(56)=>mul_re_out(1822),
            data_re_in(57)=>mul_re_out(1854),
            data_re_in(58)=>mul_re_out(1886),
            data_re_in(59)=>mul_re_out(1918),
            data_re_in(60)=>mul_re_out(1950),
            data_re_in(61)=>mul_re_out(1982),
            data_re_in(62)=>mul_re_out(2014),
            data_re_in(63)=>mul_re_out(2046),
            data_im_in(0)=>mul_im_out(30),
            data_im_in(1)=>mul_im_out(62),
            data_im_in(2)=>mul_im_out(94),
            data_im_in(3)=>mul_im_out(126),
            data_im_in(4)=>mul_im_out(158),
            data_im_in(5)=>mul_im_out(190),
            data_im_in(6)=>mul_im_out(222),
            data_im_in(7)=>mul_im_out(254),
            data_im_in(8)=>mul_im_out(286),
            data_im_in(9)=>mul_im_out(318),
            data_im_in(10)=>mul_im_out(350),
            data_im_in(11)=>mul_im_out(382),
            data_im_in(12)=>mul_im_out(414),
            data_im_in(13)=>mul_im_out(446),
            data_im_in(14)=>mul_im_out(478),
            data_im_in(15)=>mul_im_out(510),
            data_im_in(16)=>mul_im_out(542),
            data_im_in(17)=>mul_im_out(574),
            data_im_in(18)=>mul_im_out(606),
            data_im_in(19)=>mul_im_out(638),
            data_im_in(20)=>mul_im_out(670),
            data_im_in(21)=>mul_im_out(702),
            data_im_in(22)=>mul_im_out(734),
            data_im_in(23)=>mul_im_out(766),
            data_im_in(24)=>mul_im_out(798),
            data_im_in(25)=>mul_im_out(830),
            data_im_in(26)=>mul_im_out(862),
            data_im_in(27)=>mul_im_out(894),
            data_im_in(28)=>mul_im_out(926),
            data_im_in(29)=>mul_im_out(958),
            data_im_in(30)=>mul_im_out(990),
            data_im_in(31)=>mul_im_out(1022),
            data_im_in(32)=>mul_im_out(1054),
            data_im_in(33)=>mul_im_out(1086),
            data_im_in(34)=>mul_im_out(1118),
            data_im_in(35)=>mul_im_out(1150),
            data_im_in(36)=>mul_im_out(1182),
            data_im_in(37)=>mul_im_out(1214),
            data_im_in(38)=>mul_im_out(1246),
            data_im_in(39)=>mul_im_out(1278),
            data_im_in(40)=>mul_im_out(1310),
            data_im_in(41)=>mul_im_out(1342),
            data_im_in(42)=>mul_im_out(1374),
            data_im_in(43)=>mul_im_out(1406),
            data_im_in(44)=>mul_im_out(1438),
            data_im_in(45)=>mul_im_out(1470),
            data_im_in(46)=>mul_im_out(1502),
            data_im_in(47)=>mul_im_out(1534),
            data_im_in(48)=>mul_im_out(1566),
            data_im_in(49)=>mul_im_out(1598),
            data_im_in(50)=>mul_im_out(1630),
            data_im_in(51)=>mul_im_out(1662),
            data_im_in(52)=>mul_im_out(1694),
            data_im_in(53)=>mul_im_out(1726),
            data_im_in(54)=>mul_im_out(1758),
            data_im_in(55)=>mul_im_out(1790),
            data_im_in(56)=>mul_im_out(1822),
            data_im_in(57)=>mul_im_out(1854),
            data_im_in(58)=>mul_im_out(1886),
            data_im_in(59)=>mul_im_out(1918),
            data_im_in(60)=>mul_im_out(1950),
            data_im_in(61)=>mul_im_out(1982),
            data_im_in(62)=>mul_im_out(2014),
            data_im_in(63)=>mul_im_out(2046),
            data_re_out(0)=>data_re_out(30),
            data_re_out(1)=>data_re_out(62),
            data_re_out(2)=>data_re_out(94),
            data_re_out(3)=>data_re_out(126),
            data_re_out(4)=>data_re_out(158),
            data_re_out(5)=>data_re_out(190),
            data_re_out(6)=>data_re_out(222),
            data_re_out(7)=>data_re_out(254),
            data_re_out(8)=>data_re_out(286),
            data_re_out(9)=>data_re_out(318),
            data_re_out(10)=>data_re_out(350),
            data_re_out(11)=>data_re_out(382),
            data_re_out(12)=>data_re_out(414),
            data_re_out(13)=>data_re_out(446),
            data_re_out(14)=>data_re_out(478),
            data_re_out(15)=>data_re_out(510),
            data_re_out(16)=>data_re_out(542),
            data_re_out(17)=>data_re_out(574),
            data_re_out(18)=>data_re_out(606),
            data_re_out(19)=>data_re_out(638),
            data_re_out(20)=>data_re_out(670),
            data_re_out(21)=>data_re_out(702),
            data_re_out(22)=>data_re_out(734),
            data_re_out(23)=>data_re_out(766),
            data_re_out(24)=>data_re_out(798),
            data_re_out(25)=>data_re_out(830),
            data_re_out(26)=>data_re_out(862),
            data_re_out(27)=>data_re_out(894),
            data_re_out(28)=>data_re_out(926),
            data_re_out(29)=>data_re_out(958),
            data_re_out(30)=>data_re_out(990),
            data_re_out(31)=>data_re_out(1022),
            data_re_out(32)=>data_re_out(1054),
            data_re_out(33)=>data_re_out(1086),
            data_re_out(34)=>data_re_out(1118),
            data_re_out(35)=>data_re_out(1150),
            data_re_out(36)=>data_re_out(1182),
            data_re_out(37)=>data_re_out(1214),
            data_re_out(38)=>data_re_out(1246),
            data_re_out(39)=>data_re_out(1278),
            data_re_out(40)=>data_re_out(1310),
            data_re_out(41)=>data_re_out(1342),
            data_re_out(42)=>data_re_out(1374),
            data_re_out(43)=>data_re_out(1406),
            data_re_out(44)=>data_re_out(1438),
            data_re_out(45)=>data_re_out(1470),
            data_re_out(46)=>data_re_out(1502),
            data_re_out(47)=>data_re_out(1534),
            data_re_out(48)=>data_re_out(1566),
            data_re_out(49)=>data_re_out(1598),
            data_re_out(50)=>data_re_out(1630),
            data_re_out(51)=>data_re_out(1662),
            data_re_out(52)=>data_re_out(1694),
            data_re_out(53)=>data_re_out(1726),
            data_re_out(54)=>data_re_out(1758),
            data_re_out(55)=>data_re_out(1790),
            data_re_out(56)=>data_re_out(1822),
            data_re_out(57)=>data_re_out(1854),
            data_re_out(58)=>data_re_out(1886),
            data_re_out(59)=>data_re_out(1918),
            data_re_out(60)=>data_re_out(1950),
            data_re_out(61)=>data_re_out(1982),
            data_re_out(62)=>data_re_out(2014),
            data_re_out(63)=>data_re_out(2046),
            data_im_out(0)=>data_im_out(30),
            data_im_out(1)=>data_im_out(62),
            data_im_out(2)=>data_im_out(94),
            data_im_out(3)=>data_im_out(126),
            data_im_out(4)=>data_im_out(158),
            data_im_out(5)=>data_im_out(190),
            data_im_out(6)=>data_im_out(222),
            data_im_out(7)=>data_im_out(254),
            data_im_out(8)=>data_im_out(286),
            data_im_out(9)=>data_im_out(318),
            data_im_out(10)=>data_im_out(350),
            data_im_out(11)=>data_im_out(382),
            data_im_out(12)=>data_im_out(414),
            data_im_out(13)=>data_im_out(446),
            data_im_out(14)=>data_im_out(478),
            data_im_out(15)=>data_im_out(510),
            data_im_out(16)=>data_im_out(542),
            data_im_out(17)=>data_im_out(574),
            data_im_out(18)=>data_im_out(606),
            data_im_out(19)=>data_im_out(638),
            data_im_out(20)=>data_im_out(670),
            data_im_out(21)=>data_im_out(702),
            data_im_out(22)=>data_im_out(734),
            data_im_out(23)=>data_im_out(766),
            data_im_out(24)=>data_im_out(798),
            data_im_out(25)=>data_im_out(830),
            data_im_out(26)=>data_im_out(862),
            data_im_out(27)=>data_im_out(894),
            data_im_out(28)=>data_im_out(926),
            data_im_out(29)=>data_im_out(958),
            data_im_out(30)=>data_im_out(990),
            data_im_out(31)=>data_im_out(1022),
            data_im_out(32)=>data_im_out(1054),
            data_im_out(33)=>data_im_out(1086),
            data_im_out(34)=>data_im_out(1118),
            data_im_out(35)=>data_im_out(1150),
            data_im_out(36)=>data_im_out(1182),
            data_im_out(37)=>data_im_out(1214),
            data_im_out(38)=>data_im_out(1246),
            data_im_out(39)=>data_im_out(1278),
            data_im_out(40)=>data_im_out(1310),
            data_im_out(41)=>data_im_out(1342),
            data_im_out(42)=>data_im_out(1374),
            data_im_out(43)=>data_im_out(1406),
            data_im_out(44)=>data_im_out(1438),
            data_im_out(45)=>data_im_out(1470),
            data_im_out(46)=>data_im_out(1502),
            data_im_out(47)=>data_im_out(1534),
            data_im_out(48)=>data_im_out(1566),
            data_im_out(49)=>data_im_out(1598),
            data_im_out(50)=>data_im_out(1630),
            data_im_out(51)=>data_im_out(1662),
            data_im_out(52)=>data_im_out(1694),
            data_im_out(53)=>data_im_out(1726),
            data_im_out(54)=>data_im_out(1758),
            data_im_out(55)=>data_im_out(1790),
            data_im_out(56)=>data_im_out(1822),
            data_im_out(57)=>data_im_out(1854),
            data_im_out(58)=>data_im_out(1886),
            data_im_out(59)=>data_im_out(1918),
            data_im_out(60)=>data_im_out(1950),
            data_im_out(61)=>data_im_out(1982),
            data_im_out(62)=>data_im_out(2014),
            data_im_out(63)=>data_im_out(2046)
        );           

    URFFT_PT64_31 : fft_pt64
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in(0)=>mul_re_out(31),
            data_re_in(1)=>mul_re_out(63),
            data_re_in(2)=>mul_re_out(95),
            data_re_in(3)=>mul_re_out(127),
            data_re_in(4)=>mul_re_out(159),
            data_re_in(5)=>mul_re_out(191),
            data_re_in(6)=>mul_re_out(223),
            data_re_in(7)=>mul_re_out(255),
            data_re_in(8)=>mul_re_out(287),
            data_re_in(9)=>mul_re_out(319),
            data_re_in(10)=>mul_re_out(351),
            data_re_in(11)=>mul_re_out(383),
            data_re_in(12)=>mul_re_out(415),
            data_re_in(13)=>mul_re_out(447),
            data_re_in(14)=>mul_re_out(479),
            data_re_in(15)=>mul_re_out(511),
            data_re_in(16)=>mul_re_out(543),
            data_re_in(17)=>mul_re_out(575),
            data_re_in(18)=>mul_re_out(607),
            data_re_in(19)=>mul_re_out(639),
            data_re_in(20)=>mul_re_out(671),
            data_re_in(21)=>mul_re_out(703),
            data_re_in(22)=>mul_re_out(735),
            data_re_in(23)=>mul_re_out(767),
            data_re_in(24)=>mul_re_out(799),
            data_re_in(25)=>mul_re_out(831),
            data_re_in(26)=>mul_re_out(863),
            data_re_in(27)=>mul_re_out(895),
            data_re_in(28)=>mul_re_out(927),
            data_re_in(29)=>mul_re_out(959),
            data_re_in(30)=>mul_re_out(991),
            data_re_in(31)=>mul_re_out(1023),
            data_re_in(32)=>mul_re_out(1055),
            data_re_in(33)=>mul_re_out(1087),
            data_re_in(34)=>mul_re_out(1119),
            data_re_in(35)=>mul_re_out(1151),
            data_re_in(36)=>mul_re_out(1183),
            data_re_in(37)=>mul_re_out(1215),
            data_re_in(38)=>mul_re_out(1247),
            data_re_in(39)=>mul_re_out(1279),
            data_re_in(40)=>mul_re_out(1311),
            data_re_in(41)=>mul_re_out(1343),
            data_re_in(42)=>mul_re_out(1375),
            data_re_in(43)=>mul_re_out(1407),
            data_re_in(44)=>mul_re_out(1439),
            data_re_in(45)=>mul_re_out(1471),
            data_re_in(46)=>mul_re_out(1503),
            data_re_in(47)=>mul_re_out(1535),
            data_re_in(48)=>mul_re_out(1567),
            data_re_in(49)=>mul_re_out(1599),
            data_re_in(50)=>mul_re_out(1631),
            data_re_in(51)=>mul_re_out(1663),
            data_re_in(52)=>mul_re_out(1695),
            data_re_in(53)=>mul_re_out(1727),
            data_re_in(54)=>mul_re_out(1759),
            data_re_in(55)=>mul_re_out(1791),
            data_re_in(56)=>mul_re_out(1823),
            data_re_in(57)=>mul_re_out(1855),
            data_re_in(58)=>mul_re_out(1887),
            data_re_in(59)=>mul_re_out(1919),
            data_re_in(60)=>mul_re_out(1951),
            data_re_in(61)=>mul_re_out(1983),
            data_re_in(62)=>mul_re_out(2015),
            data_re_in(63)=>mul_re_out(2047),
            data_im_in(0)=>mul_im_out(31),
            data_im_in(1)=>mul_im_out(63),
            data_im_in(2)=>mul_im_out(95),
            data_im_in(3)=>mul_im_out(127),
            data_im_in(4)=>mul_im_out(159),
            data_im_in(5)=>mul_im_out(191),
            data_im_in(6)=>mul_im_out(223),
            data_im_in(7)=>mul_im_out(255),
            data_im_in(8)=>mul_im_out(287),
            data_im_in(9)=>mul_im_out(319),
            data_im_in(10)=>mul_im_out(351),
            data_im_in(11)=>mul_im_out(383),
            data_im_in(12)=>mul_im_out(415),
            data_im_in(13)=>mul_im_out(447),
            data_im_in(14)=>mul_im_out(479),
            data_im_in(15)=>mul_im_out(511),
            data_im_in(16)=>mul_im_out(543),
            data_im_in(17)=>mul_im_out(575),
            data_im_in(18)=>mul_im_out(607),
            data_im_in(19)=>mul_im_out(639),
            data_im_in(20)=>mul_im_out(671),
            data_im_in(21)=>mul_im_out(703),
            data_im_in(22)=>mul_im_out(735),
            data_im_in(23)=>mul_im_out(767),
            data_im_in(24)=>mul_im_out(799),
            data_im_in(25)=>mul_im_out(831),
            data_im_in(26)=>mul_im_out(863),
            data_im_in(27)=>mul_im_out(895),
            data_im_in(28)=>mul_im_out(927),
            data_im_in(29)=>mul_im_out(959),
            data_im_in(30)=>mul_im_out(991),
            data_im_in(31)=>mul_im_out(1023),
            data_im_in(32)=>mul_im_out(1055),
            data_im_in(33)=>mul_im_out(1087),
            data_im_in(34)=>mul_im_out(1119),
            data_im_in(35)=>mul_im_out(1151),
            data_im_in(36)=>mul_im_out(1183),
            data_im_in(37)=>mul_im_out(1215),
            data_im_in(38)=>mul_im_out(1247),
            data_im_in(39)=>mul_im_out(1279),
            data_im_in(40)=>mul_im_out(1311),
            data_im_in(41)=>mul_im_out(1343),
            data_im_in(42)=>mul_im_out(1375),
            data_im_in(43)=>mul_im_out(1407),
            data_im_in(44)=>mul_im_out(1439),
            data_im_in(45)=>mul_im_out(1471),
            data_im_in(46)=>mul_im_out(1503),
            data_im_in(47)=>mul_im_out(1535),
            data_im_in(48)=>mul_im_out(1567),
            data_im_in(49)=>mul_im_out(1599),
            data_im_in(50)=>mul_im_out(1631),
            data_im_in(51)=>mul_im_out(1663),
            data_im_in(52)=>mul_im_out(1695),
            data_im_in(53)=>mul_im_out(1727),
            data_im_in(54)=>mul_im_out(1759),
            data_im_in(55)=>mul_im_out(1791),
            data_im_in(56)=>mul_im_out(1823),
            data_im_in(57)=>mul_im_out(1855),
            data_im_in(58)=>mul_im_out(1887),
            data_im_in(59)=>mul_im_out(1919),
            data_im_in(60)=>mul_im_out(1951),
            data_im_in(61)=>mul_im_out(1983),
            data_im_in(62)=>mul_im_out(2015),
            data_im_in(63)=>mul_im_out(2047),
            data_re_out(0)=>data_re_out(31),
            data_re_out(1)=>data_re_out(63),
            data_re_out(2)=>data_re_out(95),
            data_re_out(3)=>data_re_out(127),
            data_re_out(4)=>data_re_out(159),
            data_re_out(5)=>data_re_out(191),
            data_re_out(6)=>data_re_out(223),
            data_re_out(7)=>data_re_out(255),
            data_re_out(8)=>data_re_out(287),
            data_re_out(9)=>data_re_out(319),
            data_re_out(10)=>data_re_out(351),
            data_re_out(11)=>data_re_out(383),
            data_re_out(12)=>data_re_out(415),
            data_re_out(13)=>data_re_out(447),
            data_re_out(14)=>data_re_out(479),
            data_re_out(15)=>data_re_out(511),
            data_re_out(16)=>data_re_out(543),
            data_re_out(17)=>data_re_out(575),
            data_re_out(18)=>data_re_out(607),
            data_re_out(19)=>data_re_out(639),
            data_re_out(20)=>data_re_out(671),
            data_re_out(21)=>data_re_out(703),
            data_re_out(22)=>data_re_out(735),
            data_re_out(23)=>data_re_out(767),
            data_re_out(24)=>data_re_out(799),
            data_re_out(25)=>data_re_out(831),
            data_re_out(26)=>data_re_out(863),
            data_re_out(27)=>data_re_out(895),
            data_re_out(28)=>data_re_out(927),
            data_re_out(29)=>data_re_out(959),
            data_re_out(30)=>data_re_out(991),
            data_re_out(31)=>data_re_out(1023),
            data_re_out(32)=>data_re_out(1055),
            data_re_out(33)=>data_re_out(1087),
            data_re_out(34)=>data_re_out(1119),
            data_re_out(35)=>data_re_out(1151),
            data_re_out(36)=>data_re_out(1183),
            data_re_out(37)=>data_re_out(1215),
            data_re_out(38)=>data_re_out(1247),
            data_re_out(39)=>data_re_out(1279),
            data_re_out(40)=>data_re_out(1311),
            data_re_out(41)=>data_re_out(1343),
            data_re_out(42)=>data_re_out(1375),
            data_re_out(43)=>data_re_out(1407),
            data_re_out(44)=>data_re_out(1439),
            data_re_out(45)=>data_re_out(1471),
            data_re_out(46)=>data_re_out(1503),
            data_re_out(47)=>data_re_out(1535),
            data_re_out(48)=>data_re_out(1567),
            data_re_out(49)=>data_re_out(1599),
            data_re_out(50)=>data_re_out(1631),
            data_re_out(51)=>data_re_out(1663),
            data_re_out(52)=>data_re_out(1695),
            data_re_out(53)=>data_re_out(1727),
            data_re_out(54)=>data_re_out(1759),
            data_re_out(55)=>data_re_out(1791),
            data_re_out(56)=>data_re_out(1823),
            data_re_out(57)=>data_re_out(1855),
            data_re_out(58)=>data_re_out(1887),
            data_re_out(59)=>data_re_out(1919),
            data_re_out(60)=>data_re_out(1951),
            data_re_out(61)=>data_re_out(1983),
            data_re_out(62)=>data_re_out(2015),
            data_re_out(63)=>data_re_out(2047),
            data_im_out(0)=>data_im_out(31),
            data_im_out(1)=>data_im_out(63),
            data_im_out(2)=>data_im_out(95),
            data_im_out(3)=>data_im_out(127),
            data_im_out(4)=>data_im_out(159),
            data_im_out(5)=>data_im_out(191),
            data_im_out(6)=>data_im_out(223),
            data_im_out(7)=>data_im_out(255),
            data_im_out(8)=>data_im_out(287),
            data_im_out(9)=>data_im_out(319),
            data_im_out(10)=>data_im_out(351),
            data_im_out(11)=>data_im_out(383),
            data_im_out(12)=>data_im_out(415),
            data_im_out(13)=>data_im_out(447),
            data_im_out(14)=>data_im_out(479),
            data_im_out(15)=>data_im_out(511),
            data_im_out(16)=>data_im_out(543),
            data_im_out(17)=>data_im_out(575),
            data_im_out(18)=>data_im_out(607),
            data_im_out(19)=>data_im_out(639),
            data_im_out(20)=>data_im_out(671),
            data_im_out(21)=>data_im_out(703),
            data_im_out(22)=>data_im_out(735),
            data_im_out(23)=>data_im_out(767),
            data_im_out(24)=>data_im_out(799),
            data_im_out(25)=>data_im_out(831),
            data_im_out(26)=>data_im_out(863),
            data_im_out(27)=>data_im_out(895),
            data_im_out(28)=>data_im_out(927),
            data_im_out(29)=>data_im_out(959),
            data_im_out(30)=>data_im_out(991),
            data_im_out(31)=>data_im_out(1023),
            data_im_out(32)=>data_im_out(1055),
            data_im_out(33)=>data_im_out(1087),
            data_im_out(34)=>data_im_out(1119),
            data_im_out(35)=>data_im_out(1151),
            data_im_out(36)=>data_im_out(1183),
            data_im_out(37)=>data_im_out(1215),
            data_im_out(38)=>data_im_out(1247),
            data_im_out(39)=>data_im_out(1279),
            data_im_out(40)=>data_im_out(1311),
            data_im_out(41)=>data_im_out(1343),
            data_im_out(42)=>data_im_out(1375),
            data_im_out(43)=>data_im_out(1407),
            data_im_out(44)=>data_im_out(1439),
            data_im_out(45)=>data_im_out(1471),
            data_im_out(46)=>data_im_out(1503),
            data_im_out(47)=>data_im_out(1535),
            data_im_out(48)=>data_im_out(1567),
            data_im_out(49)=>data_im_out(1599),
            data_im_out(50)=>data_im_out(1631),
            data_im_out(51)=>data_im_out(1663),
            data_im_out(52)=>data_im_out(1695),
            data_im_out(53)=>data_im_out(1727),
            data_im_out(54)=>data_im_out(1759),
            data_im_out(55)=>data_im_out(1791),
            data_im_out(56)=>data_im_out(1823),
            data_im_out(57)=>data_im_out(1855),
            data_im_out(58)=>data_im_out(1887),
            data_im_out(59)=>data_im_out(1919),
            data_im_out(60)=>data_im_out(1951),
            data_im_out(61)=>data_im_out(1983),
            data_im_out(62)=>data_im_out(2015),
            data_im_out(63)=>data_im_out(2047)
        );           


    --- multipliers
    UDELAY_0_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(0),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(0)
        );
    UDELAY_0_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(0),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(0)
        );
    USHIFTER_0_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(0),
            data_out=>mul_re_out(0)
        );
    USHIFTER_0_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(0),
            data_out=>mul_im_out(0)
        );

    UDELAY_1_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1)
        );
    UDELAY_1_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1)
        );
    USHIFTER_1_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1),
            data_out=>mul_re_out(1)
        );
    USHIFTER_1_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1),
            data_out=>mul_im_out(1)
        );

    UDELAY_2_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(2),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(2)
        );
    UDELAY_2_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(2),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(2)
        );
    USHIFTER_2_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(2),
            data_out=>mul_re_out(2)
        );
    USHIFTER_2_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(2),
            data_out=>mul_im_out(2)
        );

    UDELAY_3_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(3),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(3)
        );
    UDELAY_3_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(3),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(3)
        );
    USHIFTER_3_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(3),
            data_out=>mul_re_out(3)
        );
    USHIFTER_3_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(3),
            data_out=>mul_im_out(3)
        );

    UDELAY_4_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(4),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(4)
        );
    UDELAY_4_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(4),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(4)
        );
    USHIFTER_4_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(4),
            data_out=>mul_re_out(4)
        );
    USHIFTER_4_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(4),
            data_out=>mul_im_out(4)
        );

    UDELAY_5_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(5),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(5)
        );
    UDELAY_5_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(5),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(5)
        );
    USHIFTER_5_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(5),
            data_out=>mul_re_out(5)
        );
    USHIFTER_5_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(5),
            data_out=>mul_im_out(5)
        );

    UDELAY_6_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(6),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(6)
        );
    UDELAY_6_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(6),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(6)
        );
    USHIFTER_6_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(6),
            data_out=>mul_re_out(6)
        );
    USHIFTER_6_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(6),
            data_out=>mul_im_out(6)
        );

    UDELAY_7_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(7),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(7)
        );
    UDELAY_7_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(7),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(7)
        );
    USHIFTER_7_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(7),
            data_out=>mul_re_out(7)
        );
    USHIFTER_7_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(7),
            data_out=>mul_im_out(7)
        );

    UDELAY_8_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(8),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(8)
        );
    UDELAY_8_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(8),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(8)
        );
    USHIFTER_8_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(8),
            data_out=>mul_re_out(8)
        );
    USHIFTER_8_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(8),
            data_out=>mul_im_out(8)
        );

    UDELAY_9_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(9),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(9)
        );
    UDELAY_9_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(9),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(9)
        );
    USHIFTER_9_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(9),
            data_out=>mul_re_out(9)
        );
    USHIFTER_9_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(9),
            data_out=>mul_im_out(9)
        );

    UDELAY_10_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(10),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(10)
        );
    UDELAY_10_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(10),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(10)
        );
    USHIFTER_10_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(10),
            data_out=>mul_re_out(10)
        );
    USHIFTER_10_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(10),
            data_out=>mul_im_out(10)
        );

    UDELAY_11_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(11),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(11)
        );
    UDELAY_11_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(11),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(11)
        );
    USHIFTER_11_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(11),
            data_out=>mul_re_out(11)
        );
    USHIFTER_11_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(11),
            data_out=>mul_im_out(11)
        );

    UDELAY_12_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(12),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(12)
        );
    UDELAY_12_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(12),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(12)
        );
    USHIFTER_12_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(12),
            data_out=>mul_re_out(12)
        );
    USHIFTER_12_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(12),
            data_out=>mul_im_out(12)
        );

    UDELAY_13_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(13),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(13)
        );
    UDELAY_13_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(13),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(13)
        );
    USHIFTER_13_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(13),
            data_out=>mul_re_out(13)
        );
    USHIFTER_13_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(13),
            data_out=>mul_im_out(13)
        );

    UDELAY_14_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(14),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(14)
        );
    UDELAY_14_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(14),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(14)
        );
    USHIFTER_14_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(14),
            data_out=>mul_re_out(14)
        );
    USHIFTER_14_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(14),
            data_out=>mul_im_out(14)
        );

    UDELAY_15_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(15),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(15)
        );
    UDELAY_15_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(15),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(15)
        );
    USHIFTER_15_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(15),
            data_out=>mul_re_out(15)
        );
    USHIFTER_15_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(15),
            data_out=>mul_im_out(15)
        );

    UDELAY_16_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(16),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(16)
        );
    UDELAY_16_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(16),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(16)
        );
    USHIFTER_16_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(16),
            data_out=>mul_re_out(16)
        );
    USHIFTER_16_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(16),
            data_out=>mul_im_out(16)
        );

    UDELAY_17_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(17),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(17)
        );
    UDELAY_17_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(17),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(17)
        );
    USHIFTER_17_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(17),
            data_out=>mul_re_out(17)
        );
    USHIFTER_17_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(17),
            data_out=>mul_im_out(17)
        );

    UDELAY_18_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(18),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(18)
        );
    UDELAY_18_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(18),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(18)
        );
    USHIFTER_18_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(18),
            data_out=>mul_re_out(18)
        );
    USHIFTER_18_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(18),
            data_out=>mul_im_out(18)
        );

    UDELAY_19_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(19),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(19)
        );
    UDELAY_19_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(19),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(19)
        );
    USHIFTER_19_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(19),
            data_out=>mul_re_out(19)
        );
    USHIFTER_19_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(19),
            data_out=>mul_im_out(19)
        );

    UDELAY_20_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(20),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(20)
        );
    UDELAY_20_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(20),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(20)
        );
    USHIFTER_20_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(20),
            data_out=>mul_re_out(20)
        );
    USHIFTER_20_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(20),
            data_out=>mul_im_out(20)
        );

    UDELAY_21_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(21),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(21)
        );
    UDELAY_21_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(21),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(21)
        );
    USHIFTER_21_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(21),
            data_out=>mul_re_out(21)
        );
    USHIFTER_21_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(21),
            data_out=>mul_im_out(21)
        );

    UDELAY_22_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(22),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(22)
        );
    UDELAY_22_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(22),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(22)
        );
    USHIFTER_22_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(22),
            data_out=>mul_re_out(22)
        );
    USHIFTER_22_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(22),
            data_out=>mul_im_out(22)
        );

    UDELAY_23_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(23),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(23)
        );
    UDELAY_23_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(23),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(23)
        );
    USHIFTER_23_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(23),
            data_out=>mul_re_out(23)
        );
    USHIFTER_23_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(23),
            data_out=>mul_im_out(23)
        );

    UDELAY_24_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(24),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(24)
        );
    UDELAY_24_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(24),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(24)
        );
    USHIFTER_24_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(24),
            data_out=>mul_re_out(24)
        );
    USHIFTER_24_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(24),
            data_out=>mul_im_out(24)
        );

    UDELAY_25_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(25),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(25)
        );
    UDELAY_25_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(25),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(25)
        );
    USHIFTER_25_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(25),
            data_out=>mul_re_out(25)
        );
    USHIFTER_25_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(25),
            data_out=>mul_im_out(25)
        );

    UDELAY_26_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(26),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(26)
        );
    UDELAY_26_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(26),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(26)
        );
    USHIFTER_26_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(26),
            data_out=>mul_re_out(26)
        );
    USHIFTER_26_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(26),
            data_out=>mul_im_out(26)
        );

    UDELAY_27_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(27),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(27)
        );
    UDELAY_27_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(27),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(27)
        );
    USHIFTER_27_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(27),
            data_out=>mul_re_out(27)
        );
    USHIFTER_27_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(27),
            data_out=>mul_im_out(27)
        );

    UDELAY_28_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(28),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(28)
        );
    UDELAY_28_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(28),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(28)
        );
    USHIFTER_28_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(28),
            data_out=>mul_re_out(28)
        );
    USHIFTER_28_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(28),
            data_out=>mul_im_out(28)
        );

    UDELAY_29_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(29),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(29)
        );
    UDELAY_29_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(29),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(29)
        );
    USHIFTER_29_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(29),
            data_out=>mul_re_out(29)
        );
    USHIFTER_29_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(29),
            data_out=>mul_im_out(29)
        );

    UDELAY_30_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(30),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(30)
        );
    UDELAY_30_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(30),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(30)
        );
    USHIFTER_30_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(30),
            data_out=>mul_re_out(30)
        );
    USHIFTER_30_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(30),
            data_out=>mul_im_out(30)
        );

    UDELAY_31_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(31),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(31)
        );
    UDELAY_31_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(31),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(31)
        );
    USHIFTER_31_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(31),
            data_out=>mul_re_out(31)
        );
    USHIFTER_31_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(31),
            data_out=>mul_im_out(31)
        );

    UDELAY_32_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(32),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(32)
        );
    UDELAY_32_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(32),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(32)
        );
    USHIFTER_32_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(32),
            data_out=>mul_re_out(32)
        );
    USHIFTER_32_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(32),
            data_out=>mul_im_out(32)
        );

    UMUL_33 : complex_multiplier
    generic map(
            re_multiplicator=>16383, --- 0.999938964844 + j-0.0030517578125
            im_multiplicator=>-50
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(33),
            data_im_in=>first_stage_im_out(33),
            product_re_out=>mul_re_out(33),
            product_im_out=>mul_im_out(33)
        );

    UMUL_34 : complex_multiplier
    generic map(
            re_multiplicator=>16383, --- 0.999938964844 + j-0.006103515625
            im_multiplicator=>-100
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(34),
            data_im_in=>first_stage_im_out(34),
            product_re_out=>mul_re_out(34),
            product_im_out=>mul_im_out(34)
        );

    UMUL_35 : complex_multiplier
    generic map(
            re_multiplicator=>16383, --- 0.999938964844 + j-0.0091552734375
            im_multiplicator=>-150
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(35),
            data_im_in=>first_stage_im_out(35),
            product_re_out=>mul_re_out(35),
            product_im_out=>mul_im_out(35)
        );

    UMUL_36 : complex_multiplier
    generic map(
            re_multiplicator=>16382, --- 0.999877929688 + j-0.0122680664062
            im_multiplicator=>-201
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(36),
            data_im_in=>first_stage_im_out(36),
            product_re_out=>mul_re_out(36),
            product_im_out=>mul_im_out(36)
        );

    UMUL_37 : complex_multiplier
    generic map(
            re_multiplicator=>16382, --- 0.999877929688 + j-0.0153198242188
            im_multiplicator=>-251
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(37),
            data_im_in=>first_stage_im_out(37),
            product_re_out=>mul_re_out(37),
            product_im_out=>mul_im_out(37)
        );

    UMUL_38 : complex_multiplier
    generic map(
            re_multiplicator=>16381, --- 0.999816894531 + j-0.0183715820312
            im_multiplicator=>-301
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(38),
            data_im_in=>first_stage_im_out(38),
            product_re_out=>mul_re_out(38),
            product_im_out=>mul_im_out(38)
        );

    UMUL_39 : complex_multiplier
    generic map(
            re_multiplicator=>16380, --- 0.999755859375 + j-0.0214233398438
            im_multiplicator=>-351
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(39),
            data_im_in=>first_stage_im_out(39),
            product_re_out=>mul_re_out(39),
            product_im_out=>mul_im_out(39)
        );

    UMUL_40 : complex_multiplier
    generic map(
            re_multiplicator=>16379, --- 0.999694824219 + j-0.0245361328125
            im_multiplicator=>-402
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(40),
            data_im_in=>first_stage_im_out(40),
            product_re_out=>mul_re_out(40),
            product_im_out=>mul_im_out(40)
        );

    UMUL_41 : complex_multiplier
    generic map(
            re_multiplicator=>16377, --- 0.999572753906 + j-0.027587890625
            im_multiplicator=>-452
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(41),
            data_im_in=>first_stage_im_out(41),
            product_re_out=>mul_re_out(41),
            product_im_out=>mul_im_out(41)
        );

    UMUL_42 : complex_multiplier
    generic map(
            re_multiplicator=>16376, --- 0.99951171875 + j-0.0306396484375
            im_multiplicator=>-502
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(42),
            data_im_in=>first_stage_im_out(42),
            product_re_out=>mul_re_out(42),
            product_im_out=>mul_im_out(42)
        );

    UMUL_43 : complex_multiplier
    generic map(
            re_multiplicator=>16374, --- 0.999389648438 + j-0.03369140625
            im_multiplicator=>-552
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(43),
            data_im_in=>first_stage_im_out(43),
            product_re_out=>mul_re_out(43),
            product_im_out=>mul_im_out(43)
        );

    UMUL_44 : complex_multiplier
    generic map(
            re_multiplicator=>16372, --- 0.999267578125 + j-0.0368041992188
            im_multiplicator=>-603
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(44),
            data_im_in=>first_stage_im_out(44),
            product_re_out=>mul_re_out(44),
            product_im_out=>mul_im_out(44)
        );

    UMUL_45 : complex_multiplier
    generic map(
            re_multiplicator=>16370, --- 0.999145507812 + j-0.0398559570312
            im_multiplicator=>-653
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(45),
            data_im_in=>first_stage_im_out(45),
            product_re_out=>mul_re_out(45),
            product_im_out=>mul_im_out(45)
        );

    UMUL_46 : complex_multiplier
    generic map(
            re_multiplicator=>16368, --- 0.9990234375 + j-0.0429077148438
            im_multiplicator=>-703
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(46),
            data_im_in=>first_stage_im_out(46),
            product_re_out=>mul_re_out(46),
            product_im_out=>mul_im_out(46)
        );

    UMUL_47 : complex_multiplier
    generic map(
            re_multiplicator=>16366, --- 0.998901367188 + j-0.0459594726562
            im_multiplicator=>-753
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(47),
            data_im_in=>first_stage_im_out(47),
            product_re_out=>mul_re_out(47),
            product_im_out=>mul_im_out(47)
        );

    UMUL_48 : complex_multiplier
    generic map(
            re_multiplicator=>16364, --- 0.998779296875 + j-0.0490112304688
            im_multiplicator=>-803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(48),
            data_im_in=>first_stage_im_out(48),
            product_re_out=>mul_re_out(48),
            product_im_out=>mul_im_out(48)
        );

    UMUL_49 : complex_multiplier
    generic map(
            re_multiplicator=>16361, --- 0.998596191406 + j-0.0521240234375
            im_multiplicator=>-854
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(49),
            data_im_in=>first_stage_im_out(49),
            product_re_out=>mul_re_out(49),
            product_im_out=>mul_im_out(49)
        );

    UMUL_50 : complex_multiplier
    generic map(
            re_multiplicator=>16359, --- 0.998474121094 + j-0.05517578125
            im_multiplicator=>-904
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(50),
            data_im_in=>first_stage_im_out(50),
            product_re_out=>mul_re_out(50),
            product_im_out=>mul_im_out(50)
        );

    UMUL_51 : complex_multiplier
    generic map(
            re_multiplicator=>16356, --- 0.998291015625 + j-0.0582275390625
            im_multiplicator=>-954
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(51),
            data_im_in=>first_stage_im_out(51),
            product_re_out=>mul_re_out(51),
            product_im_out=>mul_im_out(51)
        );

    UMUL_52 : complex_multiplier
    generic map(
            re_multiplicator=>16353, --- 0.998107910156 + j-0.061279296875
            im_multiplicator=>-1004
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(52),
            data_im_in=>first_stage_im_out(52),
            product_re_out=>mul_re_out(52),
            product_im_out=>mul_im_out(52)
        );

    UMUL_53 : complex_multiplier
    generic map(
            re_multiplicator=>16350, --- 0.997924804688 + j-0.0643310546875
            im_multiplicator=>-1054
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(53),
            data_im_in=>first_stage_im_out(53),
            product_re_out=>mul_re_out(53),
            product_im_out=>mul_im_out(53)
        );

    UMUL_54 : complex_multiplier
    generic map(
            re_multiplicator=>16346, --- 0.997680664062 + j-0.0674438476562
            im_multiplicator=>-1105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(54),
            data_im_in=>first_stage_im_out(54),
            product_re_out=>mul_re_out(54),
            product_im_out=>mul_im_out(54)
        );

    UMUL_55 : complex_multiplier
    generic map(
            re_multiplicator=>16343, --- 0.997497558594 + j-0.0704956054688
            im_multiplicator=>-1155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(55),
            data_im_in=>first_stage_im_out(55),
            product_re_out=>mul_re_out(55),
            product_im_out=>mul_im_out(55)
        );

    UMUL_56 : complex_multiplier
    generic map(
            re_multiplicator=>16339, --- 0.997253417969 + j-0.0735473632812
            im_multiplicator=>-1205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(56),
            data_im_in=>first_stage_im_out(56),
            product_re_out=>mul_re_out(56),
            product_im_out=>mul_im_out(56)
        );

    UMUL_57 : complex_multiplier
    generic map(
            re_multiplicator=>16335, --- 0.997009277344 + j-0.0765991210938
            im_multiplicator=>-1255
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(57),
            data_im_in=>first_stage_im_out(57),
            product_re_out=>mul_re_out(57),
            product_im_out=>mul_im_out(57)
        );

    UMUL_58 : complex_multiplier
    generic map(
            re_multiplicator=>16331, --- 0.996765136719 + j-0.0796508789062
            im_multiplicator=>-1305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(58),
            data_im_in=>first_stage_im_out(58),
            product_re_out=>mul_re_out(58),
            product_im_out=>mul_im_out(58)
        );

    UMUL_59 : complex_multiplier
    generic map(
            re_multiplicator=>16327, --- 0.996520996094 + j-0.0827026367188
            im_multiplicator=>-1355
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(59),
            data_im_in=>first_stage_im_out(59),
            product_re_out=>mul_re_out(59),
            product_im_out=>mul_im_out(59)
        );

    UMUL_60 : complex_multiplier
    generic map(
            re_multiplicator=>16323, --- 0.996276855469 + j-0.0857543945312
            im_multiplicator=>-1405
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(60),
            data_im_in=>first_stage_im_out(60),
            product_re_out=>mul_re_out(60),
            product_im_out=>mul_im_out(60)
        );

    UMUL_61 : complex_multiplier
    generic map(
            re_multiplicator=>16319, --- 0.996032714844 + j-0.0888061523438
            im_multiplicator=>-1455
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(61),
            data_im_in=>first_stage_im_out(61),
            product_re_out=>mul_re_out(61),
            product_im_out=>mul_im_out(61)
        );

    UMUL_62 : complex_multiplier
    generic map(
            re_multiplicator=>16314, --- 0.995727539062 + j-0.0918579101562
            im_multiplicator=>-1505
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(62),
            data_im_in=>first_stage_im_out(62),
            product_re_out=>mul_re_out(62),
            product_im_out=>mul_im_out(62)
        );

    UMUL_63 : complex_multiplier
    generic map(
            re_multiplicator=>16309, --- 0.995422363281 + j-0.0949096679688
            im_multiplicator=>-1555
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(63),
            data_im_in=>first_stage_im_out(63),
            product_re_out=>mul_re_out(63),
            product_im_out=>mul_im_out(63)
        );

    UDELAY_64_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(64),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(64)
        );
    UDELAY_64_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(64),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(64)
        );
    USHIFTER_64_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(64),
            data_out=>mul_re_out(64)
        );
    USHIFTER_64_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(64),
            data_out=>mul_im_out(64)
        );

    UMUL_65 : complex_multiplier
    generic map(
            re_multiplicator=>16383, --- 0.999938964844 + j-0.006103515625
            im_multiplicator=>-100
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(65),
            data_im_in=>first_stage_im_out(65),
            product_re_out=>mul_re_out(65),
            product_im_out=>mul_im_out(65)
        );

    UMUL_66 : complex_multiplier
    generic map(
            re_multiplicator=>16382, --- 0.999877929688 + j-0.0122680664062
            im_multiplicator=>-201
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(66),
            data_im_in=>first_stage_im_out(66),
            product_re_out=>mul_re_out(66),
            product_im_out=>mul_im_out(66)
        );

    UMUL_67 : complex_multiplier
    generic map(
            re_multiplicator=>16381, --- 0.999816894531 + j-0.0183715820312
            im_multiplicator=>-301
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(67),
            data_im_in=>first_stage_im_out(67),
            product_re_out=>mul_re_out(67),
            product_im_out=>mul_im_out(67)
        );

    UMUL_68 : complex_multiplier
    generic map(
            re_multiplicator=>16379, --- 0.999694824219 + j-0.0245361328125
            im_multiplicator=>-402
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(68),
            data_im_in=>first_stage_im_out(68),
            product_re_out=>mul_re_out(68),
            product_im_out=>mul_im_out(68)
        );

    UMUL_69 : complex_multiplier
    generic map(
            re_multiplicator=>16376, --- 0.99951171875 + j-0.0306396484375
            im_multiplicator=>-502
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(69),
            data_im_in=>first_stage_im_out(69),
            product_re_out=>mul_re_out(69),
            product_im_out=>mul_im_out(69)
        );

    UMUL_70 : complex_multiplier
    generic map(
            re_multiplicator=>16372, --- 0.999267578125 + j-0.0368041992188
            im_multiplicator=>-603
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(70),
            data_im_in=>first_stage_im_out(70),
            product_re_out=>mul_re_out(70),
            product_im_out=>mul_im_out(70)
        );

    UMUL_71 : complex_multiplier
    generic map(
            re_multiplicator=>16368, --- 0.9990234375 + j-0.0429077148438
            im_multiplicator=>-703
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(71),
            data_im_in=>first_stage_im_out(71),
            product_re_out=>mul_re_out(71),
            product_im_out=>mul_im_out(71)
        );

    UMUL_72 : complex_multiplier
    generic map(
            re_multiplicator=>16364, --- 0.998779296875 + j-0.0490112304688
            im_multiplicator=>-803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(72),
            data_im_in=>first_stage_im_out(72),
            product_re_out=>mul_re_out(72),
            product_im_out=>mul_im_out(72)
        );

    UMUL_73 : complex_multiplier
    generic map(
            re_multiplicator=>16359, --- 0.998474121094 + j-0.05517578125
            im_multiplicator=>-904
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(73),
            data_im_in=>first_stage_im_out(73),
            product_re_out=>mul_re_out(73),
            product_im_out=>mul_im_out(73)
        );

    UMUL_74 : complex_multiplier
    generic map(
            re_multiplicator=>16353, --- 0.998107910156 + j-0.061279296875
            im_multiplicator=>-1004
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(74),
            data_im_in=>first_stage_im_out(74),
            product_re_out=>mul_re_out(74),
            product_im_out=>mul_im_out(74)
        );

    UMUL_75 : complex_multiplier
    generic map(
            re_multiplicator=>16346, --- 0.997680664062 + j-0.0674438476562
            im_multiplicator=>-1105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(75),
            data_im_in=>first_stage_im_out(75),
            product_re_out=>mul_re_out(75),
            product_im_out=>mul_im_out(75)
        );

    UMUL_76 : complex_multiplier
    generic map(
            re_multiplicator=>16339, --- 0.997253417969 + j-0.0735473632812
            im_multiplicator=>-1205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(76),
            data_im_in=>first_stage_im_out(76),
            product_re_out=>mul_re_out(76),
            product_im_out=>mul_im_out(76)
        );

    UMUL_77 : complex_multiplier
    generic map(
            re_multiplicator=>16331, --- 0.996765136719 + j-0.0796508789062
            im_multiplicator=>-1305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(77),
            data_im_in=>first_stage_im_out(77),
            product_re_out=>mul_re_out(77),
            product_im_out=>mul_im_out(77)
        );

    UMUL_78 : complex_multiplier
    generic map(
            re_multiplicator=>16323, --- 0.996276855469 + j-0.0857543945312
            im_multiplicator=>-1405
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(78),
            data_im_in=>first_stage_im_out(78),
            product_re_out=>mul_re_out(78),
            product_im_out=>mul_im_out(78)
        );

    UMUL_79 : complex_multiplier
    generic map(
            re_multiplicator=>16314, --- 0.995727539062 + j-0.0918579101562
            im_multiplicator=>-1505
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(79),
            data_im_in=>first_stage_im_out(79),
            product_re_out=>mul_re_out(79),
            product_im_out=>mul_im_out(79)
        );

    UMUL_80 : complex_multiplier
    generic map(
            re_multiplicator=>16305, --- 0.995178222656 + j-0.0979614257812
            im_multiplicator=>-1605
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(80),
            data_im_in=>first_stage_im_out(80),
            product_re_out=>mul_re_out(80),
            product_im_out=>mul_im_out(80)
        );

    UMUL_81 : complex_multiplier
    generic map(
            re_multiplicator=>16294, --- 0.994506835938 + j-0.104064941406
            im_multiplicator=>-1705
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(81),
            data_im_in=>first_stage_im_out(81),
            product_re_out=>mul_re_out(81),
            product_im_out=>mul_im_out(81)
        );

    UMUL_82 : complex_multiplier
    generic map(
            re_multiplicator=>16284, --- 0.993896484375 + j-0.110168457031
            im_multiplicator=>-1805
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(82),
            data_im_in=>first_stage_im_out(82),
            product_re_out=>mul_re_out(82),
            product_im_out=>mul_im_out(82)
        );

    UMUL_83 : complex_multiplier
    generic map(
            re_multiplicator=>16272, --- 0.9931640625 + j-0.116271972656
            im_multiplicator=>-1905
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(83),
            data_im_in=>first_stage_im_out(83),
            product_re_out=>mul_re_out(83),
            product_im_out=>mul_im_out(83)
        );

    UMUL_84 : complex_multiplier
    generic map(
            re_multiplicator=>16260, --- 0.992431640625 + j-0.122375488281
            im_multiplicator=>-2005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(84),
            data_im_in=>first_stage_im_out(84),
            product_re_out=>mul_re_out(84),
            product_im_out=>mul_im_out(84)
        );

    UMUL_85 : complex_multiplier
    generic map(
            re_multiplicator=>16248, --- 0.99169921875 + j-0.128479003906
            im_multiplicator=>-2105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(85),
            data_im_in=>first_stage_im_out(85),
            product_re_out=>mul_re_out(85),
            product_im_out=>mul_im_out(85)
        );

    UMUL_86 : complex_multiplier
    generic map(
            re_multiplicator=>16234, --- 0.990844726562 + j-0.134521484375
            im_multiplicator=>-2204
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(86),
            data_im_in=>first_stage_im_out(86),
            product_re_out=>mul_re_out(86),
            product_im_out=>mul_im_out(86)
        );

    UMUL_87 : complex_multiplier
    generic map(
            re_multiplicator=>16221, --- 0.990051269531 + j-0.140625
            im_multiplicator=>-2304
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(87),
            data_im_in=>first_stage_im_out(87),
            product_re_out=>mul_re_out(87),
            product_im_out=>mul_im_out(87)
        );

    UMUL_88 : complex_multiplier
    generic map(
            re_multiplicator=>16206, --- 0.989135742188 + j-0.146728515625
            im_multiplicator=>-2404
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(88),
            data_im_in=>first_stage_im_out(88),
            product_re_out=>mul_re_out(88),
            product_im_out=>mul_im_out(88)
        );

    UMUL_89 : complex_multiplier
    generic map(
            re_multiplicator=>16191, --- 0.988220214844 + j-0.152770996094
            im_multiplicator=>-2503
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(89),
            data_im_in=>first_stage_im_out(89),
            product_re_out=>mul_re_out(89),
            product_im_out=>mul_im_out(89)
        );

    UMUL_90 : complex_multiplier
    generic map(
            re_multiplicator=>16175, --- 0.987243652344 + j-0.158813476562
            im_multiplicator=>-2602
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(90),
            data_im_in=>first_stage_im_out(90),
            product_re_out=>mul_re_out(90),
            product_im_out=>mul_im_out(90)
        );

    UMUL_91 : complex_multiplier
    generic map(
            re_multiplicator=>16159, --- 0.986267089844 + j-0.164855957031
            im_multiplicator=>-2701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(91),
            data_im_in=>first_stage_im_out(91),
            product_re_out=>mul_re_out(91),
            product_im_out=>mul_im_out(91)
        );

    UMUL_92 : complex_multiplier
    generic map(
            re_multiplicator=>16142, --- 0.985229492188 + j-0.170959472656
            im_multiplicator=>-2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(92),
            data_im_in=>first_stage_im_out(92),
            product_re_out=>mul_re_out(92),
            product_im_out=>mul_im_out(92)
        );

    UMUL_93 : complex_multiplier
    generic map(
            re_multiplicator=>16125, --- 0.984191894531 + j-0.177001953125
            im_multiplicator=>-2900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(93),
            data_im_in=>first_stage_im_out(93),
            product_re_out=>mul_re_out(93),
            product_im_out=>mul_im_out(93)
        );

    UMUL_94 : complex_multiplier
    generic map(
            re_multiplicator=>16107, --- 0.983093261719 + j-0.182983398438
            im_multiplicator=>-2998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(94),
            data_im_in=>first_stage_im_out(94),
            product_re_out=>mul_re_out(94),
            product_im_out=>mul_im_out(94)
        );

    UMUL_95 : complex_multiplier
    generic map(
            re_multiplicator=>16088, --- 0.98193359375 + j-0.189025878906
            im_multiplicator=>-3097
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(95),
            data_im_in=>first_stage_im_out(95),
            product_re_out=>mul_re_out(95),
            product_im_out=>mul_im_out(95)
        );

    UDELAY_96_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(96),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(96)
        );
    UDELAY_96_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(96),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(96)
        );
    USHIFTER_96_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(96),
            data_out=>mul_re_out(96)
        );
    USHIFTER_96_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(96),
            data_out=>mul_im_out(96)
        );

    UMUL_97 : complex_multiplier
    generic map(
            re_multiplicator=>16383, --- 0.999938964844 + j-0.0091552734375
            im_multiplicator=>-150
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(97),
            data_im_in=>first_stage_im_out(97),
            product_re_out=>mul_re_out(97),
            product_im_out=>mul_im_out(97)
        );

    UMUL_98 : complex_multiplier
    generic map(
            re_multiplicator=>16381, --- 0.999816894531 + j-0.0183715820312
            im_multiplicator=>-301
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(98),
            data_im_in=>first_stage_im_out(98),
            product_re_out=>mul_re_out(98),
            product_im_out=>mul_im_out(98)
        );

    UMUL_99 : complex_multiplier
    generic map(
            re_multiplicator=>16377, --- 0.999572753906 + j-0.027587890625
            im_multiplicator=>-452
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(99),
            data_im_in=>first_stage_im_out(99),
            product_re_out=>mul_re_out(99),
            product_im_out=>mul_im_out(99)
        );

    UMUL_100 : complex_multiplier
    generic map(
            re_multiplicator=>16372, --- 0.999267578125 + j-0.0368041992188
            im_multiplicator=>-603
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(100),
            data_im_in=>first_stage_im_out(100),
            product_re_out=>mul_re_out(100),
            product_im_out=>mul_im_out(100)
        );

    UMUL_101 : complex_multiplier
    generic map(
            re_multiplicator=>16366, --- 0.998901367188 + j-0.0459594726562
            im_multiplicator=>-753
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(101),
            data_im_in=>first_stage_im_out(101),
            product_re_out=>mul_re_out(101),
            product_im_out=>mul_im_out(101)
        );

    UMUL_102 : complex_multiplier
    generic map(
            re_multiplicator=>16359, --- 0.998474121094 + j-0.05517578125
            im_multiplicator=>-904
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(102),
            data_im_in=>first_stage_im_out(102),
            product_re_out=>mul_re_out(102),
            product_im_out=>mul_im_out(102)
        );

    UMUL_103 : complex_multiplier
    generic map(
            re_multiplicator=>16350, --- 0.997924804688 + j-0.0643310546875
            im_multiplicator=>-1054
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(103),
            data_im_in=>first_stage_im_out(103),
            product_re_out=>mul_re_out(103),
            product_im_out=>mul_im_out(103)
        );

    UMUL_104 : complex_multiplier
    generic map(
            re_multiplicator=>16339, --- 0.997253417969 + j-0.0735473632812
            im_multiplicator=>-1205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(104),
            data_im_in=>first_stage_im_out(104),
            product_re_out=>mul_re_out(104),
            product_im_out=>mul_im_out(104)
        );

    UMUL_105 : complex_multiplier
    generic map(
            re_multiplicator=>16327, --- 0.996520996094 + j-0.0827026367188
            im_multiplicator=>-1355
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(105),
            data_im_in=>first_stage_im_out(105),
            product_re_out=>mul_re_out(105),
            product_im_out=>mul_im_out(105)
        );

    UMUL_106 : complex_multiplier
    generic map(
            re_multiplicator=>16314, --- 0.995727539062 + j-0.0918579101562
            im_multiplicator=>-1505
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(106),
            data_im_in=>first_stage_im_out(106),
            product_re_out=>mul_re_out(106),
            product_im_out=>mul_im_out(106)
        );

    UMUL_107 : complex_multiplier
    generic map(
            re_multiplicator=>16300, --- 0.994873046875 + j-0.101013183594
            im_multiplicator=>-1655
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(107),
            data_im_in=>first_stage_im_out(107),
            product_re_out=>mul_re_out(107),
            product_im_out=>mul_im_out(107)
        );

    UMUL_108 : complex_multiplier
    generic map(
            re_multiplicator=>16284, --- 0.993896484375 + j-0.110168457031
            im_multiplicator=>-1805
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(108),
            data_im_in=>first_stage_im_out(108),
            product_re_out=>mul_re_out(108),
            product_im_out=>mul_im_out(108)
        );

    UMUL_109 : complex_multiplier
    generic map(
            re_multiplicator=>16266, --- 0.992797851562 + j-0.119323730469
            im_multiplicator=>-1955
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(109),
            data_im_in=>first_stage_im_out(109),
            product_re_out=>mul_re_out(109),
            product_im_out=>mul_im_out(109)
        );

    UMUL_110 : complex_multiplier
    generic map(
            re_multiplicator=>16248, --- 0.99169921875 + j-0.128479003906
            im_multiplicator=>-2105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(110),
            data_im_in=>first_stage_im_out(110),
            product_re_out=>mul_re_out(110),
            product_im_out=>mul_im_out(110)
        );

    UMUL_111 : complex_multiplier
    generic map(
            re_multiplicator=>16228, --- 0.990478515625 + j-0.137573242188
            im_multiplicator=>-2254
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(111),
            data_im_in=>first_stage_im_out(111),
            product_re_out=>mul_re_out(111),
            product_im_out=>mul_im_out(111)
        );

    UMUL_112 : complex_multiplier
    generic map(
            re_multiplicator=>16206, --- 0.989135742188 + j-0.146728515625
            im_multiplicator=>-2404
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(112),
            data_im_in=>first_stage_im_out(112),
            product_re_out=>mul_re_out(112),
            product_im_out=>mul_im_out(112)
        );

    UMUL_113 : complex_multiplier
    generic map(
            re_multiplicator=>16183, --- 0.987731933594 + j-0.155822753906
            im_multiplicator=>-2553
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(113),
            data_im_in=>first_stage_im_out(113),
            product_re_out=>mul_re_out(113),
            product_im_out=>mul_im_out(113)
        );

    UMUL_114 : complex_multiplier
    generic map(
            re_multiplicator=>16159, --- 0.986267089844 + j-0.164855957031
            im_multiplicator=>-2701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(114),
            data_im_in=>first_stage_im_out(114),
            product_re_out=>mul_re_out(114),
            product_im_out=>mul_im_out(114)
        );

    UMUL_115 : complex_multiplier
    generic map(
            re_multiplicator=>16134, --- 0.984741210938 + j-0.173950195312
            im_multiplicator=>-2850
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(115),
            data_im_in=>first_stage_im_out(115),
            product_re_out=>mul_re_out(115),
            product_im_out=>mul_im_out(115)
        );

    UMUL_116 : complex_multiplier
    generic map(
            re_multiplicator=>16107, --- 0.983093261719 + j-0.182983398438
            im_multiplicator=>-2998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(116),
            data_im_in=>first_stage_im_out(116),
            product_re_out=>mul_re_out(116),
            product_im_out=>mul_im_out(116)
        );

    UMUL_117 : complex_multiplier
    generic map(
            re_multiplicator=>16078, --- 0.981323242188 + j-0.192077636719
            im_multiplicator=>-3147
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(117),
            data_im_in=>first_stage_im_out(117),
            product_re_out=>mul_re_out(117),
            product_im_out=>mul_im_out(117)
        );

    UMUL_118 : complex_multiplier
    generic map(
            re_multiplicator=>16049, --- 0.979553222656 + j-0.201049804688
            im_multiplicator=>-3294
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(118),
            data_im_in=>first_stage_im_out(118),
            product_re_out=>mul_re_out(118),
            product_im_out=>mul_im_out(118)
        );

    UMUL_119 : complex_multiplier
    generic map(
            re_multiplicator=>16018, --- 0.977661132812 + j-0.210083007812
            im_multiplicator=>-3442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(119),
            data_im_in=>first_stage_im_out(119),
            product_re_out=>mul_re_out(119),
            product_im_out=>mul_im_out(119)
        );

    UMUL_120 : complex_multiplier
    generic map(
            re_multiplicator=>15985, --- 0.975646972656 + j-0.219055175781
            im_multiplicator=>-3589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(120),
            data_im_in=>first_stage_im_out(120),
            product_re_out=>mul_re_out(120),
            product_im_out=>mul_im_out(120)
        );

    UMUL_121 : complex_multiplier
    generic map(
            re_multiplicator=>15952, --- 0.9736328125 + j-0.22802734375
            im_multiplicator=>-3736
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(121),
            data_im_in=>first_stage_im_out(121),
            product_re_out=>mul_re_out(121),
            product_im_out=>mul_im_out(121)
        );

    UMUL_122 : complex_multiplier
    generic map(
            re_multiplicator=>15917, --- 0.971496582031 + j-0.236999511719
            im_multiplicator=>-3883
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(122),
            data_im_in=>first_stage_im_out(122),
            product_re_out=>mul_re_out(122),
            product_im_out=>mul_im_out(122)
        );

    UMUL_123 : complex_multiplier
    generic map(
            re_multiplicator=>15880, --- 0.96923828125 + j-0.245910644531
            im_multiplicator=>-4029
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(123),
            data_im_in=>first_stage_im_out(123),
            product_re_out=>mul_re_out(123),
            product_im_out=>mul_im_out(123)
        );

    UMUL_124 : complex_multiplier
    generic map(
            re_multiplicator=>15842, --- 0.966918945312 + j-0.254821777344
            im_multiplicator=>-4175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(124),
            data_im_in=>first_stage_im_out(124),
            product_re_out=>mul_re_out(124),
            product_im_out=>mul_im_out(124)
        );

    UMUL_125 : complex_multiplier
    generic map(
            re_multiplicator=>15803, --- 0.964538574219 + j-0.263732910156
            im_multiplicator=>-4321
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(125),
            data_im_in=>first_stage_im_out(125),
            product_re_out=>mul_re_out(125),
            product_im_out=>mul_im_out(125)
        );

    UMUL_126 : complex_multiplier
    generic map(
            re_multiplicator=>15763, --- 0.962097167969 + j-0.272583007812
            im_multiplicator=>-4466
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(126),
            data_im_in=>first_stage_im_out(126),
            product_re_out=>mul_re_out(126),
            product_im_out=>mul_im_out(126)
        );

    UMUL_127 : complex_multiplier
    generic map(
            re_multiplicator=>15721, --- 0.959533691406 + j-0.281433105469
            im_multiplicator=>-4611
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(127),
            data_im_in=>first_stage_im_out(127),
            product_re_out=>mul_re_out(127),
            product_im_out=>mul_im_out(127)
        );

    UDELAY_128_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(128),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(128)
        );
    UDELAY_128_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(128),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(128)
        );
    USHIFTER_128_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(128),
            data_out=>mul_re_out(128)
        );
    USHIFTER_128_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(128),
            data_out=>mul_im_out(128)
        );

    UMUL_129 : complex_multiplier
    generic map(
            re_multiplicator=>16382, --- 0.999877929688 + j-0.0122680664062
            im_multiplicator=>-201
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(129),
            data_im_in=>first_stage_im_out(129),
            product_re_out=>mul_re_out(129),
            product_im_out=>mul_im_out(129)
        );

    UMUL_130 : complex_multiplier
    generic map(
            re_multiplicator=>16379, --- 0.999694824219 + j-0.0245361328125
            im_multiplicator=>-402
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(130),
            data_im_in=>first_stage_im_out(130),
            product_re_out=>mul_re_out(130),
            product_im_out=>mul_im_out(130)
        );

    UMUL_131 : complex_multiplier
    generic map(
            re_multiplicator=>16372, --- 0.999267578125 + j-0.0368041992188
            im_multiplicator=>-603
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(131),
            data_im_in=>first_stage_im_out(131),
            product_re_out=>mul_re_out(131),
            product_im_out=>mul_im_out(131)
        );

    UMUL_132 : complex_multiplier
    generic map(
            re_multiplicator=>16364, --- 0.998779296875 + j-0.0490112304688
            im_multiplicator=>-803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(132),
            data_im_in=>first_stage_im_out(132),
            product_re_out=>mul_re_out(132),
            product_im_out=>mul_im_out(132)
        );

    UMUL_133 : complex_multiplier
    generic map(
            re_multiplicator=>16353, --- 0.998107910156 + j-0.061279296875
            im_multiplicator=>-1004
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(133),
            data_im_in=>first_stage_im_out(133),
            product_re_out=>mul_re_out(133),
            product_im_out=>mul_im_out(133)
        );

    UMUL_134 : complex_multiplier
    generic map(
            re_multiplicator=>16339, --- 0.997253417969 + j-0.0735473632812
            im_multiplicator=>-1205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(134),
            data_im_in=>first_stage_im_out(134),
            product_re_out=>mul_re_out(134),
            product_im_out=>mul_im_out(134)
        );

    UMUL_135 : complex_multiplier
    generic map(
            re_multiplicator=>16323, --- 0.996276855469 + j-0.0857543945312
            im_multiplicator=>-1405
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(135),
            data_im_in=>first_stage_im_out(135),
            product_re_out=>mul_re_out(135),
            product_im_out=>mul_im_out(135)
        );

    UMUL_136 : complex_multiplier
    generic map(
            re_multiplicator=>16305, --- 0.995178222656 + j-0.0979614257812
            im_multiplicator=>-1605
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(136),
            data_im_in=>first_stage_im_out(136),
            product_re_out=>mul_re_out(136),
            product_im_out=>mul_im_out(136)
        );

    UMUL_137 : complex_multiplier
    generic map(
            re_multiplicator=>16284, --- 0.993896484375 + j-0.110168457031
            im_multiplicator=>-1805
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(137),
            data_im_in=>first_stage_im_out(137),
            product_re_out=>mul_re_out(137),
            product_im_out=>mul_im_out(137)
        );

    UMUL_138 : complex_multiplier
    generic map(
            re_multiplicator=>16260, --- 0.992431640625 + j-0.122375488281
            im_multiplicator=>-2005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(138),
            data_im_in=>first_stage_im_out(138),
            product_re_out=>mul_re_out(138),
            product_im_out=>mul_im_out(138)
        );

    UMUL_139 : complex_multiplier
    generic map(
            re_multiplicator=>16234, --- 0.990844726562 + j-0.134521484375
            im_multiplicator=>-2204
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(139),
            data_im_in=>first_stage_im_out(139),
            product_re_out=>mul_re_out(139),
            product_im_out=>mul_im_out(139)
        );

    UMUL_140 : complex_multiplier
    generic map(
            re_multiplicator=>16206, --- 0.989135742188 + j-0.146728515625
            im_multiplicator=>-2404
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(140),
            data_im_in=>first_stage_im_out(140),
            product_re_out=>mul_re_out(140),
            product_im_out=>mul_im_out(140)
        );

    UMUL_141 : complex_multiplier
    generic map(
            re_multiplicator=>16175, --- 0.987243652344 + j-0.158813476562
            im_multiplicator=>-2602
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(141),
            data_im_in=>first_stage_im_out(141),
            product_re_out=>mul_re_out(141),
            product_im_out=>mul_im_out(141)
        );

    UMUL_142 : complex_multiplier
    generic map(
            re_multiplicator=>16142, --- 0.985229492188 + j-0.170959472656
            im_multiplicator=>-2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(142),
            data_im_in=>first_stage_im_out(142),
            product_re_out=>mul_re_out(142),
            product_im_out=>mul_im_out(142)
        );

    UMUL_143 : complex_multiplier
    generic map(
            re_multiplicator=>16107, --- 0.983093261719 + j-0.182983398438
            im_multiplicator=>-2998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(143),
            data_im_in=>first_stage_im_out(143),
            product_re_out=>mul_re_out(143),
            product_im_out=>mul_im_out(143)
        );

    UMUL_144 : complex_multiplier
    generic map(
            re_multiplicator=>16069, --- 0.980773925781 + j-0.195068359375
            im_multiplicator=>-3196
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(144),
            data_im_in=>first_stage_im_out(144),
            product_re_out=>mul_re_out(144),
            product_im_out=>mul_im_out(144)
        );

    UMUL_145 : complex_multiplier
    generic map(
            re_multiplicator=>16028, --- 0.978271484375 + j-0.207092285156
            im_multiplicator=>-3393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(145),
            data_im_in=>first_stage_im_out(145),
            product_re_out=>mul_re_out(145),
            product_im_out=>mul_im_out(145)
        );

    UMUL_146 : complex_multiplier
    generic map(
            re_multiplicator=>15985, --- 0.975646972656 + j-0.219055175781
            im_multiplicator=>-3589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(146),
            data_im_in=>first_stage_im_out(146),
            product_re_out=>mul_re_out(146),
            product_im_out=>mul_im_out(146)
        );

    UMUL_147 : complex_multiplier
    generic map(
            re_multiplicator=>15940, --- 0.972900390625 + j-0.231018066406
            im_multiplicator=>-3785
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(147),
            data_im_in=>first_stage_im_out(147),
            product_re_out=>mul_re_out(147),
            product_im_out=>mul_im_out(147)
        );

    UMUL_148 : complex_multiplier
    generic map(
            re_multiplicator=>15892, --- 0.969970703125 + j-0.242919921875
            im_multiplicator=>-3980
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(148),
            data_im_in=>first_stage_im_out(148),
            product_re_out=>mul_re_out(148),
            product_im_out=>mul_im_out(148)
        );

    UMUL_149 : complex_multiplier
    generic map(
            re_multiplicator=>15842, --- 0.966918945312 + j-0.254821777344
            im_multiplicator=>-4175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(149),
            data_im_in=>first_stage_im_out(149),
            product_re_out=>mul_re_out(149),
            product_im_out=>mul_im_out(149)
        );

    UMUL_150 : complex_multiplier
    generic map(
            re_multiplicator=>15790, --- 0.963745117188 + j-0.266662597656
            im_multiplicator=>-4369
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(150),
            data_im_in=>first_stage_im_out(150),
            product_re_out=>mul_re_out(150),
            product_im_out=>mul_im_out(150)
        );

    UMUL_151 : complex_multiplier
    generic map(
            re_multiplicator=>15735, --- 0.960388183594 + j-0.278503417969
            im_multiplicator=>-4563
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(151),
            data_im_in=>first_stage_im_out(151),
            product_re_out=>mul_re_out(151),
            product_im_out=>mul_im_out(151)
        );

    UMUL_152 : complex_multiplier
    generic map(
            re_multiplicator=>15678, --- 0.956909179688 + j-0.290283203125
            im_multiplicator=>-4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(152),
            data_im_in=>first_stage_im_out(152),
            product_re_out=>mul_re_out(152),
            product_im_out=>mul_im_out(152)
        );

    UMUL_153 : complex_multiplier
    generic map(
            re_multiplicator=>15618, --- 0.953247070312 + j-0.302001953125
            im_multiplicator=>-4948
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(153),
            data_im_in=>first_stage_im_out(153),
            product_re_out=>mul_re_out(153),
            product_im_out=>mul_im_out(153)
        );

    UMUL_154 : complex_multiplier
    generic map(
            re_multiplicator=>15557, --- 0.949523925781 + j-0.313659667969
            im_multiplicator=>-5139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(154),
            data_im_in=>first_stage_im_out(154),
            product_re_out=>mul_re_out(154),
            product_im_out=>mul_im_out(154)
        );

    UMUL_155 : complex_multiplier
    generic map(
            re_multiplicator=>15492, --- 0.945556640625 + j-0.325256347656
            im_multiplicator=>-5329
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(155),
            data_im_in=>first_stage_im_out(155),
            product_re_out=>mul_re_out(155),
            product_im_out=>mul_im_out(155)
        );

    UMUL_156 : complex_multiplier
    generic map(
            re_multiplicator=>15426, --- 0.941528320312 + j-0.336853027344
            im_multiplicator=>-5519
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(156),
            data_im_in=>first_stage_im_out(156),
            product_re_out=>mul_re_out(156),
            product_im_out=>mul_im_out(156)
        );

    UMUL_157 : complex_multiplier
    generic map(
            re_multiplicator=>15357, --- 0.937316894531 + j-0.348388671875
            im_multiplicator=>-5708
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(157),
            data_im_in=>first_stage_im_out(157),
            product_re_out=>mul_re_out(157),
            product_im_out=>mul_im_out(157)
        );

    UMUL_158 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(158),
            data_im_in=>first_stage_im_out(158),
            product_re_out=>mul_re_out(158),
            product_im_out=>mul_im_out(158)
        );

    UMUL_159 : complex_multiplier
    generic map(
            re_multiplicator=>15212, --- 0.928466796875 + j-0.371276855469
            im_multiplicator=>-6083
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(159),
            data_im_in=>first_stage_im_out(159),
            product_re_out=>mul_re_out(159),
            product_im_out=>mul_im_out(159)
        );

    UDELAY_160_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(160),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(160)
        );
    UDELAY_160_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(160),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(160)
        );
    USHIFTER_160_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(160),
            data_out=>mul_re_out(160)
        );
    USHIFTER_160_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(160),
            data_out=>mul_im_out(160)
        );

    UMUL_161 : complex_multiplier
    generic map(
            re_multiplicator=>16382, --- 0.999877929688 + j-0.0153198242188
            im_multiplicator=>-251
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(161),
            data_im_in=>first_stage_im_out(161),
            product_re_out=>mul_re_out(161),
            product_im_out=>mul_im_out(161)
        );

    UMUL_162 : complex_multiplier
    generic map(
            re_multiplicator=>16376, --- 0.99951171875 + j-0.0306396484375
            im_multiplicator=>-502
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(162),
            data_im_in=>first_stage_im_out(162),
            product_re_out=>mul_re_out(162),
            product_im_out=>mul_im_out(162)
        );

    UMUL_163 : complex_multiplier
    generic map(
            re_multiplicator=>16366, --- 0.998901367188 + j-0.0459594726562
            im_multiplicator=>-753
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(163),
            data_im_in=>first_stage_im_out(163),
            product_re_out=>mul_re_out(163),
            product_im_out=>mul_im_out(163)
        );

    UMUL_164 : complex_multiplier
    generic map(
            re_multiplicator=>16353, --- 0.998107910156 + j-0.061279296875
            im_multiplicator=>-1004
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(164),
            data_im_in=>first_stage_im_out(164),
            product_re_out=>mul_re_out(164),
            product_im_out=>mul_im_out(164)
        );

    UMUL_165 : complex_multiplier
    generic map(
            re_multiplicator=>16335, --- 0.997009277344 + j-0.0765991210938
            im_multiplicator=>-1255
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(165),
            data_im_in=>first_stage_im_out(165),
            product_re_out=>mul_re_out(165),
            product_im_out=>mul_im_out(165)
        );

    UMUL_166 : complex_multiplier
    generic map(
            re_multiplicator=>16314, --- 0.995727539062 + j-0.0918579101562
            im_multiplicator=>-1505
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(166),
            data_im_in=>first_stage_im_out(166),
            product_re_out=>mul_re_out(166),
            product_im_out=>mul_im_out(166)
        );

    UMUL_167 : complex_multiplier
    generic map(
            re_multiplicator=>16289, --- 0.994201660156 + j-0.107116699219
            im_multiplicator=>-1755
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(167),
            data_im_in=>first_stage_im_out(167),
            product_re_out=>mul_re_out(167),
            product_im_out=>mul_im_out(167)
        );

    UMUL_168 : complex_multiplier
    generic map(
            re_multiplicator=>16260, --- 0.992431640625 + j-0.122375488281
            im_multiplicator=>-2005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(168),
            data_im_in=>first_stage_im_out(168),
            product_re_out=>mul_re_out(168),
            product_im_out=>mul_im_out(168)
        );

    UMUL_169 : complex_multiplier
    generic map(
            re_multiplicator=>16228, --- 0.990478515625 + j-0.137573242188
            im_multiplicator=>-2254
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(169),
            data_im_in=>first_stage_im_out(169),
            product_re_out=>mul_re_out(169),
            product_im_out=>mul_im_out(169)
        );

    UMUL_170 : complex_multiplier
    generic map(
            re_multiplicator=>16191, --- 0.988220214844 + j-0.152770996094
            im_multiplicator=>-2503
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(170),
            data_im_in=>first_stage_im_out(170),
            product_re_out=>mul_re_out(170),
            product_im_out=>mul_im_out(170)
        );

    UMUL_171 : complex_multiplier
    generic map(
            re_multiplicator=>16151, --- 0.985778808594 + j-0.167907714844
            im_multiplicator=>-2751
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(171),
            data_im_in=>first_stage_im_out(171),
            product_re_out=>mul_re_out(171),
            product_im_out=>mul_im_out(171)
        );

    UMUL_172 : complex_multiplier
    generic map(
            re_multiplicator=>16107, --- 0.983093261719 + j-0.182983398438
            im_multiplicator=>-2998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(172),
            data_im_in=>first_stage_im_out(172),
            product_re_out=>mul_re_out(172),
            product_im_out=>mul_im_out(172)
        );

    UMUL_173 : complex_multiplier
    generic map(
            re_multiplicator=>16059, --- 0.980163574219 + j-0.198059082031
            im_multiplicator=>-3245
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(173),
            data_im_in=>first_stage_im_out(173),
            product_re_out=>mul_re_out(173),
            product_im_out=>mul_im_out(173)
        );

    UMUL_174 : complex_multiplier
    generic map(
            re_multiplicator=>16007, --- 0.976989746094 + j-0.213073730469
            im_multiplicator=>-3491
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(174),
            data_im_in=>first_stage_im_out(174),
            product_re_out=>mul_re_out(174),
            product_im_out=>mul_im_out(174)
        );

    UMUL_175 : complex_multiplier
    generic map(
            re_multiplicator=>15952, --- 0.9736328125 + j-0.22802734375
            im_multiplicator=>-3736
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(175),
            data_im_in=>first_stage_im_out(175),
            product_re_out=>mul_re_out(175),
            product_im_out=>mul_im_out(175)
        );

    UMUL_176 : complex_multiplier
    generic map(
            re_multiplicator=>15892, --- 0.969970703125 + j-0.242919921875
            im_multiplicator=>-3980
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(176),
            data_im_in=>first_stage_im_out(176),
            product_re_out=>mul_re_out(176),
            product_im_out=>mul_im_out(176)
        );

    UMUL_177 : complex_multiplier
    generic map(
            re_multiplicator=>15830, --- 0.966186523438 + j-0.2578125
            im_multiplicator=>-4224
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(177),
            data_im_in=>first_stage_im_out(177),
            product_re_out=>mul_re_out(177),
            product_im_out=>mul_im_out(177)
        );

    UMUL_178 : complex_multiplier
    generic map(
            re_multiplicator=>15763, --- 0.962097167969 + j-0.272583007812
            im_multiplicator=>-4466
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(178),
            data_im_in=>first_stage_im_out(178),
            product_re_out=>mul_re_out(178),
            product_im_out=>mul_im_out(178)
        );

    UMUL_179 : complex_multiplier
    generic map(
            re_multiplicator=>15693, --- 0.957824707031 + j-0.287292480469
            im_multiplicator=>-4707
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(179),
            data_im_in=>first_stage_im_out(179),
            product_re_out=>mul_re_out(179),
            product_im_out=>mul_im_out(179)
        );

    UMUL_180 : complex_multiplier
    generic map(
            re_multiplicator=>15618, --- 0.953247070312 + j-0.302001953125
            im_multiplicator=>-4948
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(180),
            data_im_in=>first_stage_im_out(180),
            product_re_out=>mul_re_out(180),
            product_im_out=>mul_im_out(180)
        );

    UMUL_181 : complex_multiplier
    generic map(
            re_multiplicator=>15541, --- 0.948547363281 + j-0.316589355469
            im_multiplicator=>-5187
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(181),
            data_im_in=>first_stage_im_out(181),
            product_re_out=>mul_re_out(181),
            product_im_out=>mul_im_out(181)
        );

    UMUL_182 : complex_multiplier
    generic map(
            re_multiplicator=>15459, --- 0.943542480469 + j-0.3310546875
            im_multiplicator=>-5424
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(182),
            data_im_in=>first_stage_im_out(182),
            product_re_out=>mul_re_out(182),
            product_im_out=>mul_im_out(182)
        );

    UMUL_183 : complex_multiplier
    generic map(
            re_multiplicator=>15374, --- 0.938354492188 + j-0.345520019531
            im_multiplicator=>-5661
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(183),
            data_im_in=>first_stage_im_out(183),
            product_re_out=>mul_re_out(183),
            product_im_out=>mul_im_out(183)
        );

    UMUL_184 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(184),
            data_im_in=>first_stage_im_out(184),
            product_re_out=>mul_re_out(184),
            product_im_out=>mul_im_out(184)
        );

    UMUL_185 : complex_multiplier
    generic map(
            re_multiplicator=>15193, --- 0.927307128906 + j-0.374145507812
            im_multiplicator=>-6130
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(185),
            data_im_in=>first_stage_im_out(185),
            product_re_out=>mul_re_out(185),
            product_im_out=>mul_im_out(185)
        );

    UMUL_186 : complex_multiplier
    generic map(
            re_multiplicator=>15098, --- 0.921508789062 + j-0.388305664062
            im_multiplicator=>-6362
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(186),
            data_im_in=>first_stage_im_out(186),
            product_re_out=>mul_re_out(186),
            product_im_out=>mul_im_out(186)
        );

    UMUL_187 : complex_multiplier
    generic map(
            re_multiplicator=>14998, --- 0.915405273438 + j-0.402404785156
            im_multiplicator=>-6593
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(187),
            data_im_in=>first_stage_im_out(187),
            product_re_out=>mul_re_out(187),
            product_im_out=>mul_im_out(187)
        );

    UMUL_188 : complex_multiplier
    generic map(
            re_multiplicator=>14895, --- 0.909118652344 + j-0.416381835938
            im_multiplicator=>-6822
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(188),
            data_im_in=>first_stage_im_out(188),
            product_re_out=>mul_re_out(188),
            product_im_out=>mul_im_out(188)
        );

    UMUL_189 : complex_multiplier
    generic map(
            re_multiplicator=>14789, --- 0.902648925781 + j-0.430297851562
            im_multiplicator=>-7050
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(189),
            data_im_in=>first_stage_im_out(189),
            product_re_out=>mul_re_out(189),
            product_im_out=>mul_im_out(189)
        );

    UMUL_190 : complex_multiplier
    generic map(
            re_multiplicator=>14679, --- 0.895935058594 + j-0.444091796875
            im_multiplicator=>-7276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(190),
            data_im_in=>first_stage_im_out(190),
            product_re_out=>mul_re_out(190),
            product_im_out=>mul_im_out(190)
        );

    UMUL_191 : complex_multiplier
    generic map(
            re_multiplicator=>14566, --- 0.889038085938 + j-0.457763671875
            im_multiplicator=>-7500
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(191),
            data_im_in=>first_stage_im_out(191),
            product_re_out=>mul_re_out(191),
            product_im_out=>mul_im_out(191)
        );

    UDELAY_192_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(192),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(192)
        );
    UDELAY_192_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(192),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(192)
        );
    USHIFTER_192_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(192),
            data_out=>mul_re_out(192)
        );
    USHIFTER_192_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(192),
            data_out=>mul_im_out(192)
        );

    UMUL_193 : complex_multiplier
    generic map(
            re_multiplicator=>16381, --- 0.999816894531 + j-0.0183715820312
            im_multiplicator=>-301
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(193),
            data_im_in=>first_stage_im_out(193),
            product_re_out=>mul_re_out(193),
            product_im_out=>mul_im_out(193)
        );

    UMUL_194 : complex_multiplier
    generic map(
            re_multiplicator=>16372, --- 0.999267578125 + j-0.0368041992188
            im_multiplicator=>-603
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(194),
            data_im_in=>first_stage_im_out(194),
            product_re_out=>mul_re_out(194),
            product_im_out=>mul_im_out(194)
        );

    UMUL_195 : complex_multiplier
    generic map(
            re_multiplicator=>16359, --- 0.998474121094 + j-0.05517578125
            im_multiplicator=>-904
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(195),
            data_im_in=>first_stage_im_out(195),
            product_re_out=>mul_re_out(195),
            product_im_out=>mul_im_out(195)
        );

    UMUL_196 : complex_multiplier
    generic map(
            re_multiplicator=>16339, --- 0.997253417969 + j-0.0735473632812
            im_multiplicator=>-1205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(196),
            data_im_in=>first_stage_im_out(196),
            product_re_out=>mul_re_out(196),
            product_im_out=>mul_im_out(196)
        );

    UMUL_197 : complex_multiplier
    generic map(
            re_multiplicator=>16314, --- 0.995727539062 + j-0.0918579101562
            im_multiplicator=>-1505
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(197),
            data_im_in=>first_stage_im_out(197),
            product_re_out=>mul_re_out(197),
            product_im_out=>mul_im_out(197)
        );

    UMUL_198 : complex_multiplier
    generic map(
            re_multiplicator=>16284, --- 0.993896484375 + j-0.110168457031
            im_multiplicator=>-1805
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(198),
            data_im_in=>first_stage_im_out(198),
            product_re_out=>mul_re_out(198),
            product_im_out=>mul_im_out(198)
        );

    UMUL_199 : complex_multiplier
    generic map(
            re_multiplicator=>16248, --- 0.99169921875 + j-0.128479003906
            im_multiplicator=>-2105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(199),
            data_im_in=>first_stage_im_out(199),
            product_re_out=>mul_re_out(199),
            product_im_out=>mul_im_out(199)
        );

    UMUL_200 : complex_multiplier
    generic map(
            re_multiplicator=>16206, --- 0.989135742188 + j-0.146728515625
            im_multiplicator=>-2404
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(200),
            data_im_in=>first_stage_im_out(200),
            product_re_out=>mul_re_out(200),
            product_im_out=>mul_im_out(200)
        );

    UMUL_201 : complex_multiplier
    generic map(
            re_multiplicator=>16159, --- 0.986267089844 + j-0.164855957031
            im_multiplicator=>-2701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(201),
            data_im_in=>first_stage_im_out(201),
            product_re_out=>mul_re_out(201),
            product_im_out=>mul_im_out(201)
        );

    UMUL_202 : complex_multiplier
    generic map(
            re_multiplicator=>16107, --- 0.983093261719 + j-0.182983398438
            im_multiplicator=>-2998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(202),
            data_im_in=>first_stage_im_out(202),
            product_re_out=>mul_re_out(202),
            product_im_out=>mul_im_out(202)
        );

    UMUL_203 : complex_multiplier
    generic map(
            re_multiplicator=>16049, --- 0.979553222656 + j-0.201049804688
            im_multiplicator=>-3294
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(203),
            data_im_in=>first_stage_im_out(203),
            product_re_out=>mul_re_out(203),
            product_im_out=>mul_im_out(203)
        );

    UMUL_204 : complex_multiplier
    generic map(
            re_multiplicator=>15985, --- 0.975646972656 + j-0.219055175781
            im_multiplicator=>-3589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(204),
            data_im_in=>first_stage_im_out(204),
            product_re_out=>mul_re_out(204),
            product_im_out=>mul_im_out(204)
        );

    UMUL_205 : complex_multiplier
    generic map(
            re_multiplicator=>15917, --- 0.971496582031 + j-0.236999511719
            im_multiplicator=>-3883
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(205),
            data_im_in=>first_stage_im_out(205),
            product_re_out=>mul_re_out(205),
            product_im_out=>mul_im_out(205)
        );

    UMUL_206 : complex_multiplier
    generic map(
            re_multiplicator=>15842, --- 0.966918945312 + j-0.254821777344
            im_multiplicator=>-4175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(206),
            data_im_in=>first_stage_im_out(206),
            product_re_out=>mul_re_out(206),
            product_im_out=>mul_im_out(206)
        );

    UMUL_207 : complex_multiplier
    generic map(
            re_multiplicator=>15763, --- 0.962097167969 + j-0.272583007812
            im_multiplicator=>-4466
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(207),
            data_im_in=>first_stage_im_out(207),
            product_re_out=>mul_re_out(207),
            product_im_out=>mul_im_out(207)
        );

    UMUL_208 : complex_multiplier
    generic map(
            re_multiplicator=>15678, --- 0.956909179688 + j-0.290283203125
            im_multiplicator=>-4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(208),
            data_im_in=>first_stage_im_out(208),
            product_re_out=>mul_re_out(208),
            product_im_out=>mul_im_out(208)
        );

    UMUL_209 : complex_multiplier
    generic map(
            re_multiplicator=>15588, --- 0.951416015625 + j-0.307800292969
            im_multiplicator=>-5043
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(209),
            data_im_in=>first_stage_im_out(209),
            product_re_out=>mul_re_out(209),
            product_im_out=>mul_im_out(209)
        );

    UMUL_210 : complex_multiplier
    generic map(
            re_multiplicator=>15492, --- 0.945556640625 + j-0.325256347656
            im_multiplicator=>-5329
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(210),
            data_im_in=>first_stage_im_out(210),
            product_re_out=>mul_re_out(210),
            product_im_out=>mul_im_out(210)
        );

    UMUL_211 : complex_multiplier
    generic map(
            re_multiplicator=>15392, --- 0.939453125 + j-0.342651367188
            im_multiplicator=>-5614
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(211),
            data_im_in=>first_stage_im_out(211),
            product_re_out=>mul_re_out(211),
            product_im_out=>mul_im_out(211)
        );

    UMUL_212 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(212),
            data_im_in=>first_stage_im_out(212),
            product_re_out=>mul_re_out(212),
            product_im_out=>mul_im_out(212)
        );

    UMUL_213 : complex_multiplier
    generic map(
            re_multiplicator=>15175, --- 0.926208496094 + j-0.376953125
            im_multiplicator=>-6176
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(213),
            data_im_in=>first_stage_im_out(213),
            product_re_out=>mul_re_out(213),
            product_im_out=>mul_im_out(213)
        );

    UMUL_214 : complex_multiplier
    generic map(
            re_multiplicator=>15058, --- 0.919067382812 + j-0.393981933594
            im_multiplicator=>-6455
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(214),
            data_im_in=>first_stage_im_out(214),
            product_re_out=>mul_re_out(214),
            product_im_out=>mul_im_out(214)
        );

    UMUL_215 : complex_multiplier
    generic map(
            re_multiplicator=>14937, --- 0.911682128906 + j-0.410827636719
            im_multiplicator=>-6731
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(215),
            data_im_in=>first_stage_im_out(215),
            product_re_out=>mul_re_out(215),
            product_im_out=>mul_im_out(215)
        );

    UMUL_216 : complex_multiplier
    generic map(
            re_multiplicator=>14810, --- 0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(216),
            data_im_in=>first_stage_im_out(216),
            product_re_out=>mul_re_out(216),
            product_im_out=>mul_im_out(216)
        );

    UMUL_217 : complex_multiplier
    generic map(
            re_multiplicator=>14679, --- 0.895935058594 + j-0.444091796875
            im_multiplicator=>-7276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(217),
            data_im_in=>first_stage_im_out(217),
            product_re_out=>mul_re_out(217),
            product_im_out=>mul_im_out(217)
        );

    UMUL_218 : complex_multiplier
    generic map(
            re_multiplicator=>14543, --- 0.887634277344 + j-0.460510253906
            im_multiplicator=>-7545
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(218),
            data_im_in=>first_stage_im_out(218),
            product_re_out=>mul_re_out(218),
            product_im_out=>mul_im_out(218)
        );

    UMUL_219 : complex_multiplier
    generic map(
            re_multiplicator=>14401, --- 0.878967285156 + j-0.476745605469
            im_multiplicator=>-7811
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(219),
            data_im_in=>first_stage_im_out(219),
            product_re_out=>mul_re_out(219),
            product_im_out=>mul_im_out(219)
        );

    UMUL_220 : complex_multiplier
    generic map(
            re_multiplicator=>14255, --- 0.870056152344 + j-0.492858886719
            im_multiplicator=>-8075
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(220),
            data_im_in=>first_stage_im_out(220),
            product_re_out=>mul_re_out(220),
            product_im_out=>mul_im_out(220)
        );

    UMUL_221 : complex_multiplier
    generic map(
            re_multiplicator=>14104, --- 0.86083984375 + j-0.5087890625
            im_multiplicator=>-8336
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(221),
            data_im_in=>first_stage_im_out(221),
            product_re_out=>mul_re_out(221),
            product_im_out=>mul_im_out(221)
        );

    UMUL_222 : complex_multiplier
    generic map(
            re_multiplicator=>13948, --- 0.851318359375 + j-0.524536132812
            im_multiplicator=>-8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(222),
            data_im_in=>first_stage_im_out(222),
            product_re_out=>mul_re_out(222),
            product_im_out=>mul_im_out(222)
        );

    UMUL_223 : complex_multiplier
    generic map(
            re_multiplicator=>13788, --- 0.841552734375 + j-0.540161132812
            im_multiplicator=>-8850
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(223),
            data_im_in=>first_stage_im_out(223),
            product_re_out=>mul_re_out(223),
            product_im_out=>mul_im_out(223)
        );

    UDELAY_224_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(224),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(224)
        );
    UDELAY_224_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(224),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(224)
        );
    USHIFTER_224_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(224),
            data_out=>mul_re_out(224)
        );
    USHIFTER_224_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(224),
            data_out=>mul_im_out(224)
        );

    UMUL_225 : complex_multiplier
    generic map(
            re_multiplicator=>16380, --- 0.999755859375 + j-0.0214233398438
            im_multiplicator=>-351
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(225),
            data_im_in=>first_stage_im_out(225),
            product_re_out=>mul_re_out(225),
            product_im_out=>mul_im_out(225)
        );

    UMUL_226 : complex_multiplier
    generic map(
            re_multiplicator=>16368, --- 0.9990234375 + j-0.0429077148438
            im_multiplicator=>-703
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(226),
            data_im_in=>first_stage_im_out(226),
            product_re_out=>mul_re_out(226),
            product_im_out=>mul_im_out(226)
        );

    UMUL_227 : complex_multiplier
    generic map(
            re_multiplicator=>16350, --- 0.997924804688 + j-0.0643310546875
            im_multiplicator=>-1054
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(227),
            data_im_in=>first_stage_im_out(227),
            product_re_out=>mul_re_out(227),
            product_im_out=>mul_im_out(227)
        );

    UMUL_228 : complex_multiplier
    generic map(
            re_multiplicator=>16323, --- 0.996276855469 + j-0.0857543945312
            im_multiplicator=>-1405
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(228),
            data_im_in=>first_stage_im_out(228),
            product_re_out=>mul_re_out(228),
            product_im_out=>mul_im_out(228)
        );

    UMUL_229 : complex_multiplier
    generic map(
            re_multiplicator=>16289, --- 0.994201660156 + j-0.107116699219
            im_multiplicator=>-1755
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(229),
            data_im_in=>first_stage_im_out(229),
            product_re_out=>mul_re_out(229),
            product_im_out=>mul_im_out(229)
        );

    UMUL_230 : complex_multiplier
    generic map(
            re_multiplicator=>16248, --- 0.99169921875 + j-0.128479003906
            im_multiplicator=>-2105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(230),
            data_im_in=>first_stage_im_out(230),
            product_re_out=>mul_re_out(230),
            product_im_out=>mul_im_out(230)
        );

    UMUL_231 : complex_multiplier
    generic map(
            re_multiplicator=>16199, --- 0.988708496094 + j-0.149719238281
            im_multiplicator=>-2453
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(231),
            data_im_in=>first_stage_im_out(231),
            product_re_out=>mul_re_out(231),
            product_im_out=>mul_im_out(231)
        );

    UMUL_232 : complex_multiplier
    generic map(
            re_multiplicator=>16142, --- 0.985229492188 + j-0.170959472656
            im_multiplicator=>-2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(232),
            data_im_in=>first_stage_im_out(232),
            product_re_out=>mul_re_out(232),
            product_im_out=>mul_im_out(232)
        );

    UMUL_233 : complex_multiplier
    generic map(
            re_multiplicator=>16078, --- 0.981323242188 + j-0.192077636719
            im_multiplicator=>-3147
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(233),
            data_im_in=>first_stage_im_out(233),
            product_re_out=>mul_re_out(233),
            product_im_out=>mul_im_out(233)
        );

    UMUL_234 : complex_multiplier
    generic map(
            re_multiplicator=>16007, --- 0.976989746094 + j-0.213073730469
            im_multiplicator=>-3491
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(234),
            data_im_in=>first_stage_im_out(234),
            product_re_out=>mul_re_out(234),
            product_im_out=>mul_im_out(234)
        );

    UMUL_235 : complex_multiplier
    generic map(
            re_multiplicator=>15928, --- 0.97216796875 + j-0.234008789062
            im_multiplicator=>-3834
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(235),
            data_im_in=>first_stage_im_out(235),
            product_re_out=>mul_re_out(235),
            product_im_out=>mul_im_out(235)
        );

    UMUL_236 : complex_multiplier
    generic map(
            re_multiplicator=>15842, --- 0.966918945312 + j-0.254821777344
            im_multiplicator=>-4175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(236),
            data_im_in=>first_stage_im_out(236),
            product_re_out=>mul_re_out(236),
            product_im_out=>mul_im_out(236)
        );

    UMUL_237 : complex_multiplier
    generic map(
            re_multiplicator=>15749, --- 0.961242675781 + j-0.275512695312
            im_multiplicator=>-4514
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(237),
            data_im_in=>first_stage_im_out(237),
            product_re_out=>mul_re_out(237),
            product_im_out=>mul_im_out(237)
        );

    UMUL_238 : complex_multiplier
    generic map(
            re_multiplicator=>15649, --- 0.955139160156 + j-0.296142578125
            im_multiplicator=>-4852
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(238),
            data_im_in=>first_stage_im_out(238),
            product_re_out=>mul_re_out(238),
            product_im_out=>mul_im_out(238)
        );

    UMUL_239 : complex_multiplier
    generic map(
            re_multiplicator=>15541, --- 0.948547363281 + j-0.316589355469
            im_multiplicator=>-5187
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(239),
            data_im_in=>first_stage_im_out(239),
            product_re_out=>mul_re_out(239),
            product_im_out=>mul_im_out(239)
        );

    UMUL_240 : complex_multiplier
    generic map(
            re_multiplicator=>15426, --- 0.941528320312 + j-0.336853027344
            im_multiplicator=>-5519
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(240),
            data_im_in=>first_stage_im_out(240),
            product_re_out=>mul_re_out(240),
            product_im_out=>mul_im_out(240)
        );

    UMUL_241 : complex_multiplier
    generic map(
            re_multiplicator=>15304, --- 0.93408203125 + j-0.356994628906
            im_multiplicator=>-5849
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(241),
            data_im_in=>first_stage_im_out(241),
            product_re_out=>mul_re_out(241),
            product_im_out=>mul_im_out(241)
        );

    UMUL_242 : complex_multiplier
    generic map(
            re_multiplicator=>15175, --- 0.926208496094 + j-0.376953125
            im_multiplicator=>-6176
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(242),
            data_im_in=>first_stage_im_out(242),
            product_re_out=>mul_re_out(242),
            product_im_out=>mul_im_out(242)
        );

    UMUL_243 : complex_multiplier
    generic map(
            re_multiplicator=>15038, --- 0.917846679688 + j-0.396789550781
            im_multiplicator=>-6501
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(243),
            data_im_in=>first_stage_im_out(243),
            product_re_out=>mul_re_out(243),
            product_im_out=>mul_im_out(243)
        );

    UMUL_244 : complex_multiplier
    generic map(
            re_multiplicator=>14895, --- 0.909118652344 + j-0.416381835938
            im_multiplicator=>-6822
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(244),
            data_im_in=>first_stage_im_out(244),
            product_re_out=>mul_re_out(244),
            product_im_out=>mul_im_out(244)
        );

    UMUL_245 : complex_multiplier
    generic map(
            re_multiplicator=>14745, --- 0.899963378906 + j-0.435852050781
            im_multiplicator=>-7141
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(245),
            data_im_in=>first_stage_im_out(245),
            product_re_out=>mul_re_out(245),
            product_im_out=>mul_im_out(245)
        );

    UMUL_246 : complex_multiplier
    generic map(
            re_multiplicator=>14589, --- 0.890441894531 + j-0.455078125
            im_multiplicator=>-7456
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(246),
            data_im_in=>first_stage_im_out(246),
            product_re_out=>mul_re_out(246),
            product_im_out=>mul_im_out(246)
        );

    UMUL_247 : complex_multiplier
    generic map(
            re_multiplicator=>14425, --- 0.880432128906 + j-0.474060058594
            im_multiplicator=>-7767
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(247),
            data_im_in=>first_stage_im_out(247),
            product_re_out=>mul_re_out(247),
            product_im_out=>mul_im_out(247)
        );

    UMUL_248 : complex_multiplier
    generic map(
            re_multiplicator=>14255, --- 0.870056152344 + j-0.492858886719
            im_multiplicator=>-8075
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(248),
            data_im_in=>first_stage_im_out(248),
            product_re_out=>mul_re_out(248),
            product_im_out=>mul_im_out(248)
        );

    UMUL_249 : complex_multiplier
    generic map(
            re_multiplicator=>14078, --- 0.859252929688 + j-0.511413574219
            im_multiplicator=>-8379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(249),
            data_im_in=>first_stage_im_out(249),
            product_re_out=>mul_re_out(249),
            product_im_out=>mul_im_out(249)
        );

    UMUL_250 : complex_multiplier
    generic map(
            re_multiplicator=>13895, --- 0.848083496094 + j-0.52978515625
            im_multiplicator=>-8680
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(250),
            data_im_in=>first_stage_im_out(250),
            product_re_out=>mul_re_out(250),
            product_im_out=>mul_im_out(250)
        );

    UMUL_251 : complex_multiplier
    generic map(
            re_multiplicator=>13705, --- 0.836486816406 + j-0.5478515625
            im_multiplicator=>-8976
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(251),
            data_im_in=>first_stage_im_out(251),
            product_re_out=>mul_re_out(251),
            product_im_out=>mul_im_out(251)
        );

    UMUL_252 : complex_multiplier
    generic map(
            re_multiplicator=>13510, --- 0.824584960938 + j-0.565673828125
            im_multiplicator=>-9268
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(252),
            data_im_in=>first_stage_im_out(252),
            product_re_out=>mul_re_out(252),
            product_im_out=>mul_im_out(252)
        );

    UMUL_253 : complex_multiplier
    generic map(
            re_multiplicator=>13307, --- 0.812194824219 + j-0.583251953125
            im_multiplicator=>-9556
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(253),
            data_im_in=>first_stage_im_out(253),
            product_re_out=>mul_re_out(253),
            product_im_out=>mul_im_out(253)
        );

    UMUL_254 : complex_multiplier
    generic map(
            re_multiplicator=>13099, --- 0.799499511719 + j-0.6005859375
            im_multiplicator=>-9840
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(254),
            data_im_in=>first_stage_im_out(254),
            product_re_out=>mul_re_out(254),
            product_im_out=>mul_im_out(254)
        );

    UMUL_255 : complex_multiplier
    generic map(
            re_multiplicator=>12885, --- 0.786437988281 + j-0.617614746094
            im_multiplicator=>-10119
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(255),
            data_im_in=>first_stage_im_out(255),
            product_re_out=>mul_re_out(255),
            product_im_out=>mul_im_out(255)
        );

    UDELAY_256_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(256),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(256)
        );
    UDELAY_256_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(256),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(256)
        );
    USHIFTER_256_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(256),
            data_out=>mul_re_out(256)
        );
    USHIFTER_256_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(256),
            data_out=>mul_im_out(256)
        );

    UMUL_257 : complex_multiplier
    generic map(
            re_multiplicator=>16379, --- 0.999694824219 + j-0.0245361328125
            im_multiplicator=>-402
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(257),
            data_im_in=>first_stage_im_out(257),
            product_re_out=>mul_re_out(257),
            product_im_out=>mul_im_out(257)
        );

    UMUL_258 : complex_multiplier
    generic map(
            re_multiplicator=>16364, --- 0.998779296875 + j-0.0490112304688
            im_multiplicator=>-803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(258),
            data_im_in=>first_stage_im_out(258),
            product_re_out=>mul_re_out(258),
            product_im_out=>mul_im_out(258)
        );

    UMUL_259 : complex_multiplier
    generic map(
            re_multiplicator=>16339, --- 0.997253417969 + j-0.0735473632812
            im_multiplicator=>-1205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(259),
            data_im_in=>first_stage_im_out(259),
            product_re_out=>mul_re_out(259),
            product_im_out=>mul_im_out(259)
        );

    UMUL_260 : complex_multiplier
    generic map(
            re_multiplicator=>16305, --- 0.995178222656 + j-0.0979614257812
            im_multiplicator=>-1605
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(260),
            data_im_in=>first_stage_im_out(260),
            product_re_out=>mul_re_out(260),
            product_im_out=>mul_im_out(260)
        );

    UMUL_261 : complex_multiplier
    generic map(
            re_multiplicator=>16260, --- 0.992431640625 + j-0.122375488281
            im_multiplicator=>-2005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(261),
            data_im_in=>first_stage_im_out(261),
            product_re_out=>mul_re_out(261),
            product_im_out=>mul_im_out(261)
        );

    UMUL_262 : complex_multiplier
    generic map(
            re_multiplicator=>16206, --- 0.989135742188 + j-0.146728515625
            im_multiplicator=>-2404
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(262),
            data_im_in=>first_stage_im_out(262),
            product_re_out=>mul_re_out(262),
            product_im_out=>mul_im_out(262)
        );

    UMUL_263 : complex_multiplier
    generic map(
            re_multiplicator=>16142, --- 0.985229492188 + j-0.170959472656
            im_multiplicator=>-2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(263),
            data_im_in=>first_stage_im_out(263),
            product_re_out=>mul_re_out(263),
            product_im_out=>mul_im_out(263)
        );

    UMUL_264 : complex_multiplier
    generic map(
            re_multiplicator=>16069, --- 0.980773925781 + j-0.195068359375
            im_multiplicator=>-3196
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(264),
            data_im_in=>first_stage_im_out(264),
            product_re_out=>mul_re_out(264),
            product_im_out=>mul_im_out(264)
        );

    UMUL_265 : complex_multiplier
    generic map(
            re_multiplicator=>15985, --- 0.975646972656 + j-0.219055175781
            im_multiplicator=>-3589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(265),
            data_im_in=>first_stage_im_out(265),
            product_re_out=>mul_re_out(265),
            product_im_out=>mul_im_out(265)
        );

    UMUL_266 : complex_multiplier
    generic map(
            re_multiplicator=>15892, --- 0.969970703125 + j-0.242919921875
            im_multiplicator=>-3980
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(266),
            data_im_in=>first_stage_im_out(266),
            product_re_out=>mul_re_out(266),
            product_im_out=>mul_im_out(266)
        );

    UMUL_267 : complex_multiplier
    generic map(
            re_multiplicator=>15790, --- 0.963745117188 + j-0.266662597656
            im_multiplicator=>-4369
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(267),
            data_im_in=>first_stage_im_out(267),
            product_re_out=>mul_re_out(267),
            product_im_out=>mul_im_out(267)
        );

    UMUL_268 : complex_multiplier
    generic map(
            re_multiplicator=>15678, --- 0.956909179688 + j-0.290283203125
            im_multiplicator=>-4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(268),
            data_im_in=>first_stage_im_out(268),
            product_re_out=>mul_re_out(268),
            product_im_out=>mul_im_out(268)
        );

    UMUL_269 : complex_multiplier
    generic map(
            re_multiplicator=>15557, --- 0.949523925781 + j-0.313659667969
            im_multiplicator=>-5139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(269),
            data_im_in=>first_stage_im_out(269),
            product_re_out=>mul_re_out(269),
            product_im_out=>mul_im_out(269)
        );

    UMUL_270 : complex_multiplier
    generic map(
            re_multiplicator=>15426, --- 0.941528320312 + j-0.336853027344
            im_multiplicator=>-5519
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(270),
            data_im_in=>first_stage_im_out(270),
            product_re_out=>mul_re_out(270),
            product_im_out=>mul_im_out(270)
        );

    UMUL_271 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(271),
            data_im_in=>first_stage_im_out(271),
            product_re_out=>mul_re_out(271),
            product_im_out=>mul_im_out(271)
        );

    UMUL_272 : complex_multiplier
    generic map(
            re_multiplicator=>15136, --- 0.923828125 + j-0.382629394531
            im_multiplicator=>-6269
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(272),
            data_im_in=>first_stage_im_out(272),
            product_re_out=>mul_re_out(272),
            product_im_out=>mul_im_out(272)
        );

    UMUL_273 : complex_multiplier
    generic map(
            re_multiplicator=>14978, --- 0.914184570312 + j-0.405212402344
            im_multiplicator=>-6639
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(273),
            data_im_in=>first_stage_im_out(273),
            product_re_out=>mul_re_out(273),
            product_im_out=>mul_im_out(273)
        );

    UMUL_274 : complex_multiplier
    generic map(
            re_multiplicator=>14810, --- 0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(274),
            data_im_in=>first_stage_im_out(274),
            product_re_out=>mul_re_out(274),
            product_im_out=>mul_im_out(274)
        );

    UMUL_275 : complex_multiplier
    generic map(
            re_multiplicator=>14634, --- 0.893188476562 + j-0.449584960938
            im_multiplicator=>-7366
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(275),
            data_im_in=>first_stage_im_out(275),
            product_re_out=>mul_re_out(275),
            product_im_out=>mul_im_out(275)
        );

    UMUL_276 : complex_multiplier
    generic map(
            re_multiplicator=>14449, --- 0.881896972656 + j-0.471374511719
            im_multiplicator=>-7723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(276),
            data_im_in=>first_stage_im_out(276),
            product_re_out=>mul_re_out(276),
            product_im_out=>mul_im_out(276)
        );

    UMUL_277 : complex_multiplier
    generic map(
            re_multiplicator=>14255, --- 0.870056152344 + j-0.492858886719
            im_multiplicator=>-8075
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(277),
            data_im_in=>first_stage_im_out(277),
            product_re_out=>mul_re_out(277),
            product_im_out=>mul_im_out(277)
        );

    UMUL_278 : complex_multiplier
    generic map(
            re_multiplicator=>14053, --- 0.857727050781 + j-0.514099121094
            im_multiplicator=>-8423
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(278),
            data_im_in=>first_stage_im_out(278),
            product_re_out=>mul_re_out(278),
            product_im_out=>mul_im_out(278)
        );

    UMUL_279 : complex_multiplier
    generic map(
            re_multiplicator=>13842, --- 0.844848632812 + j-0.534973144531
            im_multiplicator=>-8765
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(279),
            data_im_in=>first_stage_im_out(279),
            product_re_out=>mul_re_out(279),
            product_im_out=>mul_im_out(279)
        );

    UMUL_280 : complex_multiplier
    generic map(
            re_multiplicator=>13622, --- 0.831420898438 + j-0.555541992188
            im_multiplicator=>-9102
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(280),
            data_im_in=>first_stage_im_out(280),
            product_re_out=>mul_re_out(280),
            product_im_out=>mul_im_out(280)
        );

    UMUL_281 : complex_multiplier
    generic map(
            re_multiplicator=>13395, --- 0.817565917969 + j-0.575805664062
            im_multiplicator=>-9434
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(281),
            data_im_in=>first_stage_im_out(281),
            product_re_out=>mul_re_out(281),
            product_im_out=>mul_im_out(281)
        );

    UMUL_282 : complex_multiplier
    generic map(
            re_multiplicator=>13159, --- 0.803161621094 + j-0.595642089844
            im_multiplicator=>-9759
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(282),
            data_im_in=>first_stage_im_out(282),
            product_re_out=>mul_re_out(282),
            product_im_out=>mul_im_out(282)
        );

    UMUL_283 : complex_multiplier
    generic map(
            re_multiplicator=>12916, --- 0.788330078125 + j-0.615173339844
            im_multiplicator=>-10079
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(283),
            data_im_in=>first_stage_im_out(283),
            product_re_out=>mul_re_out(283),
            product_im_out=>mul_im_out(283)
        );

    UMUL_284 : complex_multiplier
    generic map(
            re_multiplicator=>12665, --- 0.773010253906 + j-0.634338378906
            im_multiplicator=>-10393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(284),
            data_im_in=>first_stage_im_out(284),
            product_re_out=>mul_re_out(284),
            product_im_out=>mul_im_out(284)
        );

    UMUL_285 : complex_multiplier
    generic map(
            re_multiplicator=>12406, --- 0.757202148438 + j-0.653137207031
            im_multiplicator=>-10701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(285),
            data_im_in=>first_stage_im_out(285),
            product_re_out=>mul_re_out(285),
            product_im_out=>mul_im_out(285)
        );

    UMUL_286 : complex_multiplier
    generic map(
            re_multiplicator=>12139, --- 0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(286),
            data_im_in=>first_stage_im_out(286),
            product_re_out=>mul_re_out(286),
            product_im_out=>mul_im_out(286)
        );

    UMUL_287 : complex_multiplier
    generic map(
            re_multiplicator=>11866, --- 0.724243164062 + j-0.689514160156
            im_multiplicator=>-11297
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(287),
            data_im_in=>first_stage_im_out(287),
            product_re_out=>mul_re_out(287),
            product_im_out=>mul_im_out(287)
        );

    UDELAY_288_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(288),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(288)
        );
    UDELAY_288_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(288),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(288)
        );
    USHIFTER_288_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(288),
            data_out=>mul_re_out(288)
        );
    USHIFTER_288_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(288),
            data_out=>mul_im_out(288)
        );

    UMUL_289 : complex_multiplier
    generic map(
            re_multiplicator=>16377, --- 0.999572753906 + j-0.027587890625
            im_multiplicator=>-452
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(289),
            data_im_in=>first_stage_im_out(289),
            product_re_out=>mul_re_out(289),
            product_im_out=>mul_im_out(289)
        );

    UMUL_290 : complex_multiplier
    generic map(
            re_multiplicator=>16359, --- 0.998474121094 + j-0.05517578125
            im_multiplicator=>-904
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(290),
            data_im_in=>first_stage_im_out(290),
            product_re_out=>mul_re_out(290),
            product_im_out=>mul_im_out(290)
        );

    UMUL_291 : complex_multiplier
    generic map(
            re_multiplicator=>16327, --- 0.996520996094 + j-0.0827026367188
            im_multiplicator=>-1355
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(291),
            data_im_in=>first_stage_im_out(291),
            product_re_out=>mul_re_out(291),
            product_im_out=>mul_im_out(291)
        );

    UMUL_292 : complex_multiplier
    generic map(
            re_multiplicator=>16284, --- 0.993896484375 + j-0.110168457031
            im_multiplicator=>-1805
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(292),
            data_im_in=>first_stage_im_out(292),
            product_re_out=>mul_re_out(292),
            product_im_out=>mul_im_out(292)
        );

    UMUL_293 : complex_multiplier
    generic map(
            re_multiplicator=>16228, --- 0.990478515625 + j-0.137573242188
            im_multiplicator=>-2254
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(293),
            data_im_in=>first_stage_im_out(293),
            product_re_out=>mul_re_out(293),
            product_im_out=>mul_im_out(293)
        );

    UMUL_294 : complex_multiplier
    generic map(
            re_multiplicator=>16159, --- 0.986267089844 + j-0.164855957031
            im_multiplicator=>-2701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(294),
            data_im_in=>first_stage_im_out(294),
            product_re_out=>mul_re_out(294),
            product_im_out=>mul_im_out(294)
        );

    UMUL_295 : complex_multiplier
    generic map(
            re_multiplicator=>16078, --- 0.981323242188 + j-0.192077636719
            im_multiplicator=>-3147
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(295),
            data_im_in=>first_stage_im_out(295),
            product_re_out=>mul_re_out(295),
            product_im_out=>mul_im_out(295)
        );

    UMUL_296 : complex_multiplier
    generic map(
            re_multiplicator=>15985, --- 0.975646972656 + j-0.219055175781
            im_multiplicator=>-3589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(296),
            data_im_in=>first_stage_im_out(296),
            product_re_out=>mul_re_out(296),
            product_im_out=>mul_im_out(296)
        );

    UMUL_297 : complex_multiplier
    generic map(
            re_multiplicator=>15880, --- 0.96923828125 + j-0.245910644531
            im_multiplicator=>-4029
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(297),
            data_im_in=>first_stage_im_out(297),
            product_re_out=>mul_re_out(297),
            product_im_out=>mul_im_out(297)
        );

    UMUL_298 : complex_multiplier
    generic map(
            re_multiplicator=>15763, --- 0.962097167969 + j-0.272583007812
            im_multiplicator=>-4466
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(298),
            data_im_in=>first_stage_im_out(298),
            product_re_out=>mul_re_out(298),
            product_im_out=>mul_im_out(298)
        );

    UMUL_299 : complex_multiplier
    generic map(
            re_multiplicator=>15634, --- 0.954223632812 + j-0.299072265625
            im_multiplicator=>-4900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(299),
            data_im_in=>first_stage_im_out(299),
            product_re_out=>mul_re_out(299),
            product_im_out=>mul_im_out(299)
        );

    UMUL_300 : complex_multiplier
    generic map(
            re_multiplicator=>15492, --- 0.945556640625 + j-0.325256347656
            im_multiplicator=>-5329
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(300),
            data_im_in=>first_stage_im_out(300),
            product_re_out=>mul_re_out(300),
            product_im_out=>mul_im_out(300)
        );

    UMUL_301 : complex_multiplier
    generic map(
            re_multiplicator=>15339, --- 0.936218261719 + j-0.351257324219
            im_multiplicator=>-5755
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(301),
            data_im_in=>first_stage_im_out(301),
            product_re_out=>mul_re_out(301),
            product_im_out=>mul_im_out(301)
        );

    UMUL_302 : complex_multiplier
    generic map(
            re_multiplicator=>15175, --- 0.926208496094 + j-0.376953125
            im_multiplicator=>-6176
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(302),
            data_im_in=>first_stage_im_out(302),
            product_re_out=>mul_re_out(302),
            product_im_out=>mul_im_out(302)
        );

    UMUL_303 : complex_multiplier
    generic map(
            re_multiplicator=>14998, --- 0.915405273438 + j-0.402404785156
            im_multiplicator=>-6593
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(303),
            data_im_in=>first_stage_im_out(303),
            product_re_out=>mul_re_out(303),
            product_im_out=>mul_im_out(303)
        );

    UMUL_304 : complex_multiplier
    generic map(
            re_multiplicator=>14810, --- 0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(304),
            data_im_in=>first_stage_im_out(304),
            product_re_out=>mul_re_out(304),
            product_im_out=>mul_im_out(304)
        );

    UMUL_305 : complex_multiplier
    generic map(
            re_multiplicator=>14611, --- 0.891784667969 + j-0.452331542969
            im_multiplicator=>-7411
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(305),
            data_im_in=>first_stage_im_out(305),
            product_re_out=>mul_re_out(305),
            product_im_out=>mul_im_out(305)
        );

    UMUL_306 : complex_multiplier
    generic map(
            re_multiplicator=>14401, --- 0.878967285156 + j-0.476745605469
            im_multiplicator=>-7811
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(306),
            data_im_in=>first_stage_im_out(306),
            product_re_out=>mul_re_out(306),
            product_im_out=>mul_im_out(306)
        );

    UMUL_307 : complex_multiplier
    generic map(
            re_multiplicator=>14180, --- 0.865478515625 + j-0.500854492188
            im_multiplicator=>-8206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(307),
            data_im_in=>first_stage_im_out(307),
            product_re_out=>mul_re_out(307),
            product_im_out=>mul_im_out(307)
        );

    UMUL_308 : complex_multiplier
    generic map(
            re_multiplicator=>13948, --- 0.851318359375 + j-0.524536132812
            im_multiplicator=>-8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(308),
            data_im_in=>first_stage_im_out(308),
            product_re_out=>mul_re_out(308),
            product_im_out=>mul_im_out(308)
        );

    UMUL_309 : complex_multiplier
    generic map(
            re_multiplicator=>13705, --- 0.836486816406 + j-0.5478515625
            im_multiplicator=>-8976
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(309),
            data_im_in=>first_stage_im_out(309),
            product_re_out=>mul_re_out(309),
            product_im_out=>mul_im_out(309)
        );

    UMUL_310 : complex_multiplier
    generic map(
            re_multiplicator=>13452, --- 0.821044921875 + j-0.570739746094
            im_multiplicator=>-9351
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(310),
            data_im_in=>first_stage_im_out(310),
            product_re_out=>mul_re_out(310),
            product_im_out=>mul_im_out(310)
        );

    UMUL_311 : complex_multiplier
    generic map(
            re_multiplicator=>13189, --- 0.804992675781 + j-0.593200683594
            im_multiplicator=>-9719
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(311),
            data_im_in=>first_stage_im_out(311),
            product_re_out=>mul_re_out(311),
            product_im_out=>mul_im_out(311)
        );

    UMUL_312 : complex_multiplier
    generic map(
            re_multiplicator=>12916, --- 0.788330078125 + j-0.615173339844
            im_multiplicator=>-10079
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(312),
            data_im_in=>first_stage_im_out(312),
            product_re_out=>mul_re_out(312),
            product_im_out=>mul_im_out(312)
        );

    UMUL_313 : complex_multiplier
    generic map(
            re_multiplicator=>12633, --- 0.771057128906 + j-0.63671875
            im_multiplicator=>-10432
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(313),
            data_im_in=>first_stage_im_out(313),
            product_re_out=>mul_re_out(313),
            product_im_out=>mul_im_out(313)
        );

    UMUL_314 : complex_multiplier
    generic map(
            re_multiplicator=>12340, --- 0.753173828125 + j-0.657775878906
            im_multiplicator=>-10777
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(314),
            data_im_in=>first_stage_im_out(314),
            product_re_out=>mul_re_out(314),
            product_im_out=>mul_im_out(314)
        );

    UMUL_315 : complex_multiplier
    generic map(
            re_multiplicator=>12037, --- 0.734680175781 + j-0.678344726562
            im_multiplicator=>-11114
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(315),
            data_im_in=>first_stage_im_out(315),
            product_re_out=>mul_re_out(315),
            product_im_out=>mul_im_out(315)
        );

    UMUL_316 : complex_multiplier
    generic map(
            re_multiplicator=>11726, --- 0.715698242188 + j-0.698364257812
            im_multiplicator=>-11442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(316),
            data_im_in=>first_stage_im_out(316),
            product_re_out=>mul_re_out(316),
            product_im_out=>mul_im_out(316)
        );

    UMUL_317 : complex_multiplier
    generic map(
            re_multiplicator=>11406, --- 0.696166992188 + j-0.717834472656
            im_multiplicator=>-11761
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(317),
            data_im_in=>first_stage_im_out(317),
            product_re_out=>mul_re_out(317),
            product_im_out=>mul_im_out(317)
        );

    UMUL_318 : complex_multiplier
    generic map(
            re_multiplicator=>11077, --- 0.676086425781 + j-0.73681640625
            im_multiplicator=>-12072
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(318),
            data_im_in=>first_stage_im_out(318),
            product_re_out=>mul_re_out(318),
            product_im_out=>mul_im_out(318)
        );

    UMUL_319 : complex_multiplier
    generic map(
            re_multiplicator=>10739, --- 0.655456542969 + j-0.755187988281
            im_multiplicator=>-12373
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(319),
            data_im_in=>first_stage_im_out(319),
            product_re_out=>mul_re_out(319),
            product_im_out=>mul_im_out(319)
        );

    UDELAY_320_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(320),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(320)
        );
    UDELAY_320_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(320),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(320)
        );
    USHIFTER_320_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(320),
            data_out=>mul_re_out(320)
        );
    USHIFTER_320_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(320),
            data_out=>mul_im_out(320)
        );

    UMUL_321 : complex_multiplier
    generic map(
            re_multiplicator=>16376, --- 0.99951171875 + j-0.0306396484375
            im_multiplicator=>-502
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(321),
            data_im_in=>first_stage_im_out(321),
            product_re_out=>mul_re_out(321),
            product_im_out=>mul_im_out(321)
        );

    UMUL_322 : complex_multiplier
    generic map(
            re_multiplicator=>16353, --- 0.998107910156 + j-0.061279296875
            im_multiplicator=>-1004
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(322),
            data_im_in=>first_stage_im_out(322),
            product_re_out=>mul_re_out(322),
            product_im_out=>mul_im_out(322)
        );

    UMUL_323 : complex_multiplier
    generic map(
            re_multiplicator=>16314, --- 0.995727539062 + j-0.0918579101562
            im_multiplicator=>-1505
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(323),
            data_im_in=>first_stage_im_out(323),
            product_re_out=>mul_re_out(323),
            product_im_out=>mul_im_out(323)
        );

    UMUL_324 : complex_multiplier
    generic map(
            re_multiplicator=>16260, --- 0.992431640625 + j-0.122375488281
            im_multiplicator=>-2005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(324),
            data_im_in=>first_stage_im_out(324),
            product_re_out=>mul_re_out(324),
            product_im_out=>mul_im_out(324)
        );

    UMUL_325 : complex_multiplier
    generic map(
            re_multiplicator=>16191, --- 0.988220214844 + j-0.152770996094
            im_multiplicator=>-2503
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(325),
            data_im_in=>first_stage_im_out(325),
            product_re_out=>mul_re_out(325),
            product_im_out=>mul_im_out(325)
        );

    UMUL_326 : complex_multiplier
    generic map(
            re_multiplicator=>16107, --- 0.983093261719 + j-0.182983398438
            im_multiplicator=>-2998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(326),
            data_im_in=>first_stage_im_out(326),
            product_re_out=>mul_re_out(326),
            product_im_out=>mul_im_out(326)
        );

    UMUL_327 : complex_multiplier
    generic map(
            re_multiplicator=>16007, --- 0.976989746094 + j-0.213073730469
            im_multiplicator=>-3491
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(327),
            data_im_in=>first_stage_im_out(327),
            product_re_out=>mul_re_out(327),
            product_im_out=>mul_im_out(327)
        );

    UMUL_328 : complex_multiplier
    generic map(
            re_multiplicator=>15892, --- 0.969970703125 + j-0.242919921875
            im_multiplicator=>-3980
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(328),
            data_im_in=>first_stage_im_out(328),
            product_re_out=>mul_re_out(328),
            product_im_out=>mul_im_out(328)
        );

    UMUL_329 : complex_multiplier
    generic map(
            re_multiplicator=>15763, --- 0.962097167969 + j-0.272583007812
            im_multiplicator=>-4466
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(329),
            data_im_in=>first_stage_im_out(329),
            product_re_out=>mul_re_out(329),
            product_im_out=>mul_im_out(329)
        );

    UMUL_330 : complex_multiplier
    generic map(
            re_multiplicator=>15618, --- 0.953247070312 + j-0.302001953125
            im_multiplicator=>-4948
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(330),
            data_im_in=>first_stage_im_out(330),
            product_re_out=>mul_re_out(330),
            product_im_out=>mul_im_out(330)
        );

    UMUL_331 : complex_multiplier
    generic map(
            re_multiplicator=>15459, --- 0.943542480469 + j-0.3310546875
            im_multiplicator=>-5424
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(331),
            data_im_in=>first_stage_im_out(331),
            product_re_out=>mul_re_out(331),
            product_im_out=>mul_im_out(331)
        );

    UMUL_332 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(332),
            data_im_in=>first_stage_im_out(332),
            product_re_out=>mul_re_out(332),
            product_im_out=>mul_im_out(332)
        );

    UMUL_333 : complex_multiplier
    generic map(
            re_multiplicator=>15098, --- 0.921508789062 + j-0.388305664062
            im_multiplicator=>-6362
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(333),
            data_im_in=>first_stage_im_out(333),
            product_re_out=>mul_re_out(333),
            product_im_out=>mul_im_out(333)
        );

    UMUL_334 : complex_multiplier
    generic map(
            re_multiplicator=>14895, --- 0.909118652344 + j-0.416381835938
            im_multiplicator=>-6822
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(334),
            data_im_in=>first_stage_im_out(334),
            product_re_out=>mul_re_out(334),
            product_im_out=>mul_im_out(334)
        );

    UMUL_335 : complex_multiplier
    generic map(
            re_multiplicator=>14679, --- 0.895935058594 + j-0.444091796875
            im_multiplicator=>-7276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(335),
            data_im_in=>first_stage_im_out(335),
            product_re_out=>mul_re_out(335),
            product_im_out=>mul_im_out(335)
        );

    UMUL_336 : complex_multiplier
    generic map(
            re_multiplicator=>14449, --- 0.881896972656 + j-0.471374511719
            im_multiplicator=>-7723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(336),
            data_im_in=>first_stage_im_out(336),
            product_re_out=>mul_re_out(336),
            product_im_out=>mul_im_out(336)
        );

    UMUL_337 : complex_multiplier
    generic map(
            re_multiplicator=>14205, --- 0.867004394531 + j-0.498168945312
            im_multiplicator=>-8162
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(337),
            data_im_in=>first_stage_im_out(337),
            product_re_out=>mul_re_out(337),
            product_im_out=>mul_im_out(337)
        );

    UMUL_338 : complex_multiplier
    generic map(
            re_multiplicator=>13948, --- 0.851318359375 + j-0.524536132812
            im_multiplicator=>-8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(338),
            data_im_in=>first_stage_im_out(338),
            product_re_out=>mul_re_out(338),
            product_im_out=>mul_im_out(338)
        );

    UMUL_339 : complex_multiplier
    generic map(
            re_multiplicator=>13678, --- 0.834838867188 + j-0.550415039062
            im_multiplicator=>-9018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(339),
            data_im_in=>first_stage_im_out(339),
            product_re_out=>mul_re_out(339),
            product_im_out=>mul_im_out(339)
        );

    UMUL_340 : complex_multiplier
    generic map(
            re_multiplicator=>13395, --- 0.817565917969 + j-0.575805664062
            im_multiplicator=>-9434
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(340),
            data_im_in=>first_stage_im_out(340),
            product_re_out=>mul_re_out(340),
            product_im_out=>mul_im_out(340)
        );

    UMUL_341 : complex_multiplier
    generic map(
            re_multiplicator=>13099, --- 0.799499511719 + j-0.6005859375
            im_multiplicator=>-9840
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(341),
            data_im_in=>first_stage_im_out(341),
            product_re_out=>mul_re_out(341),
            product_im_out=>mul_im_out(341)
        );

    UMUL_342 : complex_multiplier
    generic map(
            re_multiplicator=>12791, --- 0.780700683594 + j-0.624816894531
            im_multiplicator=>-10237
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(342),
            data_im_in=>first_stage_im_out(342),
            product_re_out=>mul_re_out(342),
            product_im_out=>mul_im_out(342)
        );

    UMUL_343 : complex_multiplier
    generic map(
            re_multiplicator=>12471, --- 0.761169433594 + j-0.648498535156
            im_multiplicator=>-10625
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(343),
            data_im_in=>first_stage_im_out(343),
            product_re_out=>mul_re_out(343),
            product_im_out=>mul_im_out(343)
        );

    UMUL_344 : complex_multiplier
    generic map(
            re_multiplicator=>12139, --- 0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(344),
            data_im_in=>first_stage_im_out(344),
            product_re_out=>mul_re_out(344),
            product_im_out=>mul_im_out(344)
        );

    UMUL_345 : complex_multiplier
    generic map(
            re_multiplicator=>11796, --- 0.719970703125 + j-0.693969726562
            im_multiplicator=>-11370
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(345),
            data_im_in=>first_stage_im_out(345),
            product_re_out=>mul_re_out(345),
            product_im_out=>mul_im_out(345)
        );

    UMUL_346 : complex_multiplier
    generic map(
            re_multiplicator=>11442, --- 0.698364257812 + j-0.715698242188
            im_multiplicator=>-11726
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(346),
            data_im_in=>first_stage_im_out(346),
            product_re_out=>mul_re_out(346),
            product_im_out=>mul_im_out(346)
        );

    UMUL_347 : complex_multiplier
    generic map(
            re_multiplicator=>11077, --- 0.676086425781 + j-0.73681640625
            im_multiplicator=>-12072
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(347),
            data_im_in=>first_stage_im_out(347),
            product_re_out=>mul_re_out(347),
            product_im_out=>mul_im_out(347)
        );

    UMUL_348 : complex_multiplier
    generic map(
            re_multiplicator=>10701, --- 0.653137207031 + j-0.757202148438
            im_multiplicator=>-12406
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(348),
            data_im_in=>first_stage_im_out(348),
            product_re_out=>mul_re_out(348),
            product_im_out=>mul_im_out(348)
        );

    UMUL_349 : complex_multiplier
    generic map(
            re_multiplicator=>10315, --- 0.629577636719 + j-0.77685546875
            im_multiplicator=>-12728
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(349),
            data_im_in=>first_stage_im_out(349),
            product_re_out=>mul_re_out(349),
            product_im_out=>mul_im_out(349)
        );

    UMUL_350 : complex_multiplier
    generic map(
            re_multiplicator=>9920, --- 0.60546875 + j-0.795776367188
            im_multiplicator=>-13038
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(350),
            data_im_in=>first_stage_im_out(350),
            product_re_out=>mul_re_out(350),
            product_im_out=>mul_im_out(350)
        );

    UMUL_351 : complex_multiplier
    generic map(
            re_multiplicator=>9516, --- 0.580810546875 + j-0.814025878906
            im_multiplicator=>-13337
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(351),
            data_im_in=>first_stage_im_out(351),
            product_re_out=>mul_re_out(351),
            product_im_out=>mul_im_out(351)
        );

    UDELAY_352_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(352),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(352)
        );
    UDELAY_352_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(352),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(352)
        );
    USHIFTER_352_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(352),
            data_out=>mul_re_out(352)
        );
    USHIFTER_352_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(352),
            data_out=>mul_im_out(352)
        );

    UMUL_353 : complex_multiplier
    generic map(
            re_multiplicator=>16374, --- 0.999389648438 + j-0.03369140625
            im_multiplicator=>-552
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(353),
            data_im_in=>first_stage_im_out(353),
            product_re_out=>mul_re_out(353),
            product_im_out=>mul_im_out(353)
        );

    UMUL_354 : complex_multiplier
    generic map(
            re_multiplicator=>16346, --- 0.997680664062 + j-0.0674438476562
            im_multiplicator=>-1105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(354),
            data_im_in=>first_stage_im_out(354),
            product_re_out=>mul_re_out(354),
            product_im_out=>mul_im_out(354)
        );

    UMUL_355 : complex_multiplier
    generic map(
            re_multiplicator=>16300, --- 0.994873046875 + j-0.101013183594
            im_multiplicator=>-1655
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(355),
            data_im_in=>first_stage_im_out(355),
            product_re_out=>mul_re_out(355),
            product_im_out=>mul_im_out(355)
        );

    UMUL_356 : complex_multiplier
    generic map(
            re_multiplicator=>16234, --- 0.990844726562 + j-0.134521484375
            im_multiplicator=>-2204
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(356),
            data_im_in=>first_stage_im_out(356),
            product_re_out=>mul_re_out(356),
            product_im_out=>mul_im_out(356)
        );

    UMUL_357 : complex_multiplier
    generic map(
            re_multiplicator=>16151, --- 0.985778808594 + j-0.167907714844
            im_multiplicator=>-2751
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(357),
            data_im_in=>first_stage_im_out(357),
            product_re_out=>mul_re_out(357),
            product_im_out=>mul_im_out(357)
        );

    UMUL_358 : complex_multiplier
    generic map(
            re_multiplicator=>16049, --- 0.979553222656 + j-0.201049804688
            im_multiplicator=>-3294
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(358),
            data_im_in=>first_stage_im_out(358),
            product_re_out=>mul_re_out(358),
            product_im_out=>mul_im_out(358)
        );

    UMUL_359 : complex_multiplier
    generic map(
            re_multiplicator=>15928, --- 0.97216796875 + j-0.234008789062
            im_multiplicator=>-3834
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(359),
            data_im_in=>first_stage_im_out(359),
            product_re_out=>mul_re_out(359),
            product_im_out=>mul_im_out(359)
        );

    UMUL_360 : complex_multiplier
    generic map(
            re_multiplicator=>15790, --- 0.963745117188 + j-0.266662597656
            im_multiplicator=>-4369
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(360),
            data_im_in=>first_stage_im_out(360),
            product_re_out=>mul_re_out(360),
            product_im_out=>mul_im_out(360)
        );

    UMUL_361 : complex_multiplier
    generic map(
            re_multiplicator=>15634, --- 0.954223632812 + j-0.299072265625
            im_multiplicator=>-4900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(361),
            data_im_in=>first_stage_im_out(361),
            product_re_out=>mul_re_out(361),
            product_im_out=>mul_im_out(361)
        );

    UMUL_362 : complex_multiplier
    generic map(
            re_multiplicator=>15459, --- 0.943542480469 + j-0.3310546875
            im_multiplicator=>-5424
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(362),
            data_im_in=>first_stage_im_out(362),
            product_re_out=>mul_re_out(362),
            product_im_out=>mul_im_out(362)
        );

    UMUL_363 : complex_multiplier
    generic map(
            re_multiplicator=>15267, --- 0.931823730469 + j-0.362731933594
            im_multiplicator=>-5943
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(363),
            data_im_in=>first_stage_im_out(363),
            product_re_out=>mul_re_out(363),
            product_im_out=>mul_im_out(363)
        );

    UMUL_364 : complex_multiplier
    generic map(
            re_multiplicator=>15058, --- 0.919067382812 + j-0.393981933594
            im_multiplicator=>-6455
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(364),
            data_im_in=>first_stage_im_out(364),
            product_re_out=>mul_re_out(364),
            product_im_out=>mul_im_out(364)
        );

    UMUL_365 : complex_multiplier
    generic map(
            re_multiplicator=>14832, --- 0.9052734375 + j-0.424743652344
            im_multiplicator=>-6959
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(365),
            data_im_in=>first_stage_im_out(365),
            product_re_out=>mul_re_out(365),
            product_im_out=>mul_im_out(365)
        );

    UMUL_366 : complex_multiplier
    generic map(
            re_multiplicator=>14589, --- 0.890441894531 + j-0.455078125
            im_multiplicator=>-7456
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(366),
            data_im_in=>first_stage_im_out(366),
            product_re_out=>mul_re_out(366),
            product_im_out=>mul_im_out(366)
        );

    UMUL_367 : complex_multiplier
    generic map(
            re_multiplicator=>14329, --- 0.874572753906 + j-0.48486328125
            im_multiplicator=>-7944
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(367),
            data_im_in=>first_stage_im_out(367),
            product_re_out=>mul_re_out(367),
            product_im_out=>mul_im_out(367)
        );

    UMUL_368 : complex_multiplier
    generic map(
            re_multiplicator=>14053, --- 0.857727050781 + j-0.514099121094
            im_multiplicator=>-8423
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(368),
            data_im_in=>first_stage_im_out(368),
            product_re_out=>mul_re_out(368),
            product_im_out=>mul_im_out(368)
        );

    UMUL_369 : complex_multiplier
    generic map(
            re_multiplicator=>13760, --- 0.83984375 + j-0.542724609375
            im_multiplicator=>-8892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(369),
            data_im_in=>first_stage_im_out(369),
            product_re_out=>mul_re_out(369),
            product_im_out=>mul_im_out(369)
        );

    UMUL_370 : complex_multiplier
    generic map(
            re_multiplicator=>13452, --- 0.821044921875 + j-0.570739746094
            im_multiplicator=>-9351
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(370),
            data_im_in=>first_stage_im_out(370),
            product_re_out=>mul_re_out(370),
            product_im_out=>mul_im_out(370)
        );

    UMUL_371 : complex_multiplier
    generic map(
            re_multiplicator=>13129, --- 0.801330566406 + j-0.59814453125
            im_multiplicator=>-9800
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(371),
            data_im_in=>first_stage_im_out(371),
            product_re_out=>mul_re_out(371),
            product_im_out=>mul_im_out(371)
        );

    UMUL_372 : complex_multiplier
    generic map(
            re_multiplicator=>12791, --- 0.780700683594 + j-0.624816894531
            im_multiplicator=>-10237
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(372),
            data_im_in=>first_stage_im_out(372),
            product_re_out=>mul_re_out(372),
            product_im_out=>mul_im_out(372)
        );

    UMUL_373 : complex_multiplier
    generic map(
            re_multiplicator=>12438, --- 0.759155273438 + j-0.650817871094
            im_multiplicator=>-10663
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(373),
            data_im_in=>first_stage_im_out(373),
            product_re_out=>mul_re_out(373),
            product_im_out=>mul_im_out(373)
        );

    UMUL_374 : complex_multiplier
    generic map(
            re_multiplicator=>12072, --- 0.73681640625 + j-0.676086425781
            im_multiplicator=>-11077
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(374),
            data_im_in=>first_stage_im_out(374),
            product_re_out=>mul_re_out(374),
            product_im_out=>mul_im_out(374)
        );

    UMUL_375 : complex_multiplier
    generic map(
            re_multiplicator=>11691, --- 0.713562011719 + j-0.700561523438
            im_multiplicator=>-11478
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(375),
            data_im_in=>first_stage_im_out(375),
            product_re_out=>mul_re_out(375),
            product_im_out=>mul_im_out(375)
        );

    UMUL_376 : complex_multiplier
    generic map(
            re_multiplicator=>11297, --- 0.689514160156 + j-0.724243164062
            im_multiplicator=>-11866
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(376),
            data_im_in=>first_stage_im_out(376),
            product_re_out=>mul_re_out(376),
            product_im_out=>mul_im_out(376)
        );

    UMUL_377 : complex_multiplier
    generic map(
            re_multiplicator=>10890, --- 0.664672851562 + j-0.7470703125
            im_multiplicator=>-12240
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(377),
            data_im_in=>first_stage_im_out(377),
            product_re_out=>mul_re_out(377),
            product_im_out=>mul_im_out(377)
        );

    UMUL_378 : complex_multiplier
    generic map(
            re_multiplicator=>10471, --- 0.639099121094 + j-0.76904296875
            im_multiplicator=>-12600
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(378),
            data_im_in=>first_stage_im_out(378),
            product_re_out=>mul_re_out(378),
            product_im_out=>mul_im_out(378)
        );

    UMUL_379 : complex_multiplier
    generic map(
            re_multiplicator=>10040, --- 0.61279296875 + j-0.790222167969
            im_multiplicator=>-12947
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(379),
            data_im_in=>first_stage_im_out(379),
            product_re_out=>mul_re_out(379),
            product_im_out=>mul_im_out(379)
        );

    UMUL_380 : complex_multiplier
    generic map(
            re_multiplicator=>9597, --- 0.585754394531 + j-0.810424804688
            im_multiplicator=>-13278
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(380),
            data_im_in=>first_stage_im_out(380),
            product_re_out=>mul_re_out(380),
            product_im_out=>mul_im_out(380)
        );

    UMUL_381 : complex_multiplier
    generic map(
            re_multiplicator=>9144, --- 0.55810546875 + j-0.829711914062
            im_multiplicator=>-13594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(381),
            data_im_in=>first_stage_im_out(381),
            product_re_out=>mul_re_out(381),
            product_im_out=>mul_im_out(381)
        );

    UMUL_382 : complex_multiplier
    generic map(
            re_multiplicator=>8680, --- 0.52978515625 + j-0.848083496094
            im_multiplicator=>-13895
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(382),
            data_im_in=>first_stage_im_out(382),
            product_re_out=>mul_re_out(382),
            product_im_out=>mul_im_out(382)
        );

    UMUL_383 : complex_multiplier
    generic map(
            re_multiplicator=>8206, --- 0.500854492188 + j-0.865478515625
            im_multiplicator=>-14180
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(383),
            data_im_in=>first_stage_im_out(383),
            product_re_out=>mul_re_out(383),
            product_im_out=>mul_im_out(383)
        );

    UDELAY_384_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(384),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(384)
        );
    UDELAY_384_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(384),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(384)
        );
    USHIFTER_384_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(384),
            data_out=>mul_re_out(384)
        );
    USHIFTER_384_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(384),
            data_out=>mul_im_out(384)
        );

    UMUL_385 : complex_multiplier
    generic map(
            re_multiplicator=>16372, --- 0.999267578125 + j-0.0368041992188
            im_multiplicator=>-603
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(385),
            data_im_in=>first_stage_im_out(385),
            product_re_out=>mul_re_out(385),
            product_im_out=>mul_im_out(385)
        );

    UMUL_386 : complex_multiplier
    generic map(
            re_multiplicator=>16339, --- 0.997253417969 + j-0.0735473632812
            im_multiplicator=>-1205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(386),
            data_im_in=>first_stage_im_out(386),
            product_re_out=>mul_re_out(386),
            product_im_out=>mul_im_out(386)
        );

    UMUL_387 : complex_multiplier
    generic map(
            re_multiplicator=>16284, --- 0.993896484375 + j-0.110168457031
            im_multiplicator=>-1805
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(387),
            data_im_in=>first_stage_im_out(387),
            product_re_out=>mul_re_out(387),
            product_im_out=>mul_im_out(387)
        );

    UMUL_388 : complex_multiplier
    generic map(
            re_multiplicator=>16206, --- 0.989135742188 + j-0.146728515625
            im_multiplicator=>-2404
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(388),
            data_im_in=>first_stage_im_out(388),
            product_re_out=>mul_re_out(388),
            product_im_out=>mul_im_out(388)
        );

    UMUL_389 : complex_multiplier
    generic map(
            re_multiplicator=>16107, --- 0.983093261719 + j-0.182983398438
            im_multiplicator=>-2998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(389),
            data_im_in=>first_stage_im_out(389),
            product_re_out=>mul_re_out(389),
            product_im_out=>mul_im_out(389)
        );

    UMUL_390 : complex_multiplier
    generic map(
            re_multiplicator=>15985, --- 0.975646972656 + j-0.219055175781
            im_multiplicator=>-3589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(390),
            data_im_in=>first_stage_im_out(390),
            product_re_out=>mul_re_out(390),
            product_im_out=>mul_im_out(390)
        );

    UMUL_391 : complex_multiplier
    generic map(
            re_multiplicator=>15842, --- 0.966918945312 + j-0.254821777344
            im_multiplicator=>-4175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(391),
            data_im_in=>first_stage_im_out(391),
            product_re_out=>mul_re_out(391),
            product_im_out=>mul_im_out(391)
        );

    UMUL_392 : complex_multiplier
    generic map(
            re_multiplicator=>15678, --- 0.956909179688 + j-0.290283203125
            im_multiplicator=>-4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(392),
            data_im_in=>first_stage_im_out(392),
            product_re_out=>mul_re_out(392),
            product_im_out=>mul_im_out(392)
        );

    UMUL_393 : complex_multiplier
    generic map(
            re_multiplicator=>15492, --- 0.945556640625 + j-0.325256347656
            im_multiplicator=>-5329
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(393),
            data_im_in=>first_stage_im_out(393),
            product_re_out=>mul_re_out(393),
            product_im_out=>mul_im_out(393)
        );

    UMUL_394 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(394),
            data_im_in=>first_stage_im_out(394),
            product_re_out=>mul_re_out(394),
            product_im_out=>mul_im_out(394)
        );

    UMUL_395 : complex_multiplier
    generic map(
            re_multiplicator=>15058, --- 0.919067382812 + j-0.393981933594
            im_multiplicator=>-6455
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(395),
            data_im_in=>first_stage_im_out(395),
            product_re_out=>mul_re_out(395),
            product_im_out=>mul_im_out(395)
        );

    UMUL_396 : complex_multiplier
    generic map(
            re_multiplicator=>14810, --- 0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(396),
            data_im_in=>first_stage_im_out(396),
            product_re_out=>mul_re_out(396),
            product_im_out=>mul_im_out(396)
        );

    UMUL_397 : complex_multiplier
    generic map(
            re_multiplicator=>14543, --- 0.887634277344 + j-0.460510253906
            im_multiplicator=>-7545
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(397),
            data_im_in=>first_stage_im_out(397),
            product_re_out=>mul_re_out(397),
            product_im_out=>mul_im_out(397)
        );

    UMUL_398 : complex_multiplier
    generic map(
            re_multiplicator=>14255, --- 0.870056152344 + j-0.492858886719
            im_multiplicator=>-8075
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(398),
            data_im_in=>first_stage_im_out(398),
            product_re_out=>mul_re_out(398),
            product_im_out=>mul_im_out(398)
        );

    UMUL_399 : complex_multiplier
    generic map(
            re_multiplicator=>13948, --- 0.851318359375 + j-0.524536132812
            im_multiplicator=>-8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(399),
            data_im_in=>first_stage_im_out(399),
            product_re_out=>mul_re_out(399),
            product_im_out=>mul_im_out(399)
        );

    UMUL_400 : complex_multiplier
    generic map(
            re_multiplicator=>13622, --- 0.831420898438 + j-0.555541992188
            im_multiplicator=>-9102
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(400),
            data_im_in=>first_stage_im_out(400),
            product_re_out=>mul_re_out(400),
            product_im_out=>mul_im_out(400)
        );

    UMUL_401 : complex_multiplier
    generic map(
            re_multiplicator=>13278, --- 0.810424804688 + j-0.585754394531
            im_multiplicator=>-9597
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(401),
            data_im_in=>first_stage_im_out(401),
            product_re_out=>mul_re_out(401),
            product_im_out=>mul_im_out(401)
        );

    UMUL_402 : complex_multiplier
    generic map(
            re_multiplicator=>12916, --- 0.788330078125 + j-0.615173339844
            im_multiplicator=>-10079
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(402),
            data_im_in=>first_stage_im_out(402),
            product_re_out=>mul_re_out(402),
            product_im_out=>mul_im_out(402)
        );

    UMUL_403 : complex_multiplier
    generic map(
            re_multiplicator=>12536, --- 0.76513671875 + j-0.643798828125
            im_multiplicator=>-10548
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(403),
            data_im_in=>first_stage_im_out(403),
            product_re_out=>mul_re_out(403),
            product_im_out=>mul_im_out(403)
        );

    UMUL_404 : complex_multiplier
    generic map(
            re_multiplicator=>12139, --- 0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(404),
            data_im_in=>first_stage_im_out(404),
            product_re_out=>mul_re_out(404),
            product_im_out=>mul_im_out(404)
        );

    UMUL_405 : complex_multiplier
    generic map(
            re_multiplicator=>11726, --- 0.715698242188 + j-0.698364257812
            im_multiplicator=>-11442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(405),
            data_im_in=>first_stage_im_out(405),
            product_re_out=>mul_re_out(405),
            product_im_out=>mul_im_out(405)
        );

    UMUL_406 : complex_multiplier
    generic map(
            re_multiplicator=>11297, --- 0.689514160156 + j-0.724243164062
            im_multiplicator=>-11866
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(406),
            data_im_in=>first_stage_im_out(406),
            product_re_out=>mul_re_out(406),
            product_im_out=>mul_im_out(406)
        );

    UMUL_407 : complex_multiplier
    generic map(
            re_multiplicator=>10853, --- 0.662414550781 + j-0.749084472656
            im_multiplicator=>-12273
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(407),
            data_im_in=>first_stage_im_out(407),
            product_re_out=>mul_re_out(407),
            product_im_out=>mul_im_out(407)
        );

    UMUL_408 : complex_multiplier
    generic map(
            re_multiplicator=>10393, --- 0.634338378906 + j-0.773010253906
            im_multiplicator=>-12665
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(408),
            data_im_in=>first_stage_im_out(408),
            product_re_out=>mul_re_out(408),
            product_im_out=>mul_im_out(408)
        );

    UMUL_409 : complex_multiplier
    generic map(
            re_multiplicator=>9920, --- 0.60546875 + j-0.795776367188
            im_multiplicator=>-13038
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(409),
            data_im_in=>first_stage_im_out(409),
            product_re_out=>mul_re_out(409),
            product_im_out=>mul_im_out(409)
        );

    UMUL_410 : complex_multiplier
    generic map(
            re_multiplicator=>9434, --- 0.575805664062 + j-0.817565917969
            im_multiplicator=>-13395
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(410),
            data_im_in=>first_stage_im_out(410),
            product_re_out=>mul_re_out(410),
            product_im_out=>mul_im_out(410)
        );

    UMUL_411 : complex_multiplier
    generic map(
            re_multiplicator=>8934, --- 0.545288085938 + j-0.838195800781
            im_multiplicator=>-13733
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(411),
            data_im_in=>first_stage_im_out(411),
            product_re_out=>mul_re_out(411),
            product_im_out=>mul_im_out(411)
        );

    UMUL_412 : complex_multiplier
    generic map(
            re_multiplicator=>8423, --- 0.514099121094 + j-0.857727050781
            im_multiplicator=>-14053
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(412),
            data_im_in=>first_stage_im_out(412),
            product_re_out=>mul_re_out(412),
            product_im_out=>mul_im_out(412)
        );

    UMUL_413 : complex_multiplier
    generic map(
            re_multiplicator=>7900, --- 0.482177734375 + j-0.876037597656
            im_multiplicator=>-14353
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(413),
            data_im_in=>first_stage_im_out(413),
            product_re_out=>mul_re_out(413),
            product_im_out=>mul_im_out(413)
        );

    UMUL_414 : complex_multiplier
    generic map(
            re_multiplicator=>7366, --- 0.449584960938 + j-0.893188476562
            im_multiplicator=>-14634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(414),
            data_im_in=>first_stage_im_out(414),
            product_re_out=>mul_re_out(414),
            product_im_out=>mul_im_out(414)
        );

    UMUL_415 : complex_multiplier
    generic map(
            re_multiplicator=>6822, --- 0.416381835938 + j-0.909118652344
            im_multiplicator=>-14895
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(415),
            data_im_in=>first_stage_im_out(415),
            product_re_out=>mul_re_out(415),
            product_im_out=>mul_im_out(415)
        );

    UDELAY_416_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(416),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(416)
        );
    UDELAY_416_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(416),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(416)
        );
    USHIFTER_416_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(416),
            data_out=>mul_re_out(416)
        );
    USHIFTER_416_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(416),
            data_out=>mul_im_out(416)
        );

    UMUL_417 : complex_multiplier
    generic map(
            re_multiplicator=>16370, --- 0.999145507812 + j-0.0398559570312
            im_multiplicator=>-653
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(417),
            data_im_in=>first_stage_im_out(417),
            product_re_out=>mul_re_out(417),
            product_im_out=>mul_im_out(417)
        );

    UMUL_418 : complex_multiplier
    generic map(
            re_multiplicator=>16331, --- 0.996765136719 + j-0.0796508789062
            im_multiplicator=>-1305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(418),
            data_im_in=>first_stage_im_out(418),
            product_re_out=>mul_re_out(418),
            product_im_out=>mul_im_out(418)
        );

    UMUL_419 : complex_multiplier
    generic map(
            re_multiplicator=>16266, --- 0.992797851562 + j-0.119323730469
            im_multiplicator=>-1955
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(419),
            data_im_in=>first_stage_im_out(419),
            product_re_out=>mul_re_out(419),
            product_im_out=>mul_im_out(419)
        );

    UMUL_420 : complex_multiplier
    generic map(
            re_multiplicator=>16175, --- 0.987243652344 + j-0.158813476562
            im_multiplicator=>-2602
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(420),
            data_im_in=>first_stage_im_out(420),
            product_re_out=>mul_re_out(420),
            product_im_out=>mul_im_out(420)
        );

    UMUL_421 : complex_multiplier
    generic map(
            re_multiplicator=>16059, --- 0.980163574219 + j-0.198059082031
            im_multiplicator=>-3245
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(421),
            data_im_in=>first_stage_im_out(421),
            product_re_out=>mul_re_out(421),
            product_im_out=>mul_im_out(421)
        );

    UMUL_422 : complex_multiplier
    generic map(
            re_multiplicator=>15917, --- 0.971496582031 + j-0.236999511719
            im_multiplicator=>-3883
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(422),
            data_im_in=>first_stage_im_out(422),
            product_re_out=>mul_re_out(422),
            product_im_out=>mul_im_out(422)
        );

    UMUL_423 : complex_multiplier
    generic map(
            re_multiplicator=>15749, --- 0.961242675781 + j-0.275512695312
            im_multiplicator=>-4514
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(423),
            data_im_in=>first_stage_im_out(423),
            product_re_out=>mul_re_out(423),
            product_im_out=>mul_im_out(423)
        );

    UMUL_424 : complex_multiplier
    generic map(
            re_multiplicator=>15557, --- 0.949523925781 + j-0.313659667969
            im_multiplicator=>-5139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(424),
            data_im_in=>first_stage_im_out(424),
            product_re_out=>mul_re_out(424),
            product_im_out=>mul_im_out(424)
        );

    UMUL_425 : complex_multiplier
    generic map(
            re_multiplicator=>15339, --- 0.936218261719 + j-0.351257324219
            im_multiplicator=>-5755
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(425),
            data_im_in=>first_stage_im_out(425),
            product_re_out=>mul_re_out(425),
            product_im_out=>mul_im_out(425)
        );

    UMUL_426 : complex_multiplier
    generic map(
            re_multiplicator=>15098, --- 0.921508789062 + j-0.388305664062
            im_multiplicator=>-6362
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(426),
            data_im_in=>first_stage_im_out(426),
            product_re_out=>mul_re_out(426),
            product_im_out=>mul_im_out(426)
        );

    UMUL_427 : complex_multiplier
    generic map(
            re_multiplicator=>14832, --- 0.9052734375 + j-0.424743652344
            im_multiplicator=>-6959
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(427),
            data_im_in=>first_stage_im_out(427),
            product_re_out=>mul_re_out(427),
            product_im_out=>mul_im_out(427)
        );

    UMUL_428 : complex_multiplier
    generic map(
            re_multiplicator=>14543, --- 0.887634277344 + j-0.460510253906
            im_multiplicator=>-7545
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(428),
            data_im_in=>first_stage_im_out(428),
            product_re_out=>mul_re_out(428),
            product_im_out=>mul_im_out(428)
        );

    UMUL_429 : complex_multiplier
    generic map(
            re_multiplicator=>14230, --- 0.868530273438 + j-0.495544433594
            im_multiplicator=>-8119
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(429),
            data_im_in=>first_stage_im_out(429),
            product_re_out=>mul_re_out(429),
            product_im_out=>mul_im_out(429)
        );

    UMUL_430 : complex_multiplier
    generic map(
            re_multiplicator=>13895, --- 0.848083496094 + j-0.52978515625
            im_multiplicator=>-8680
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(430),
            data_im_in=>first_stage_im_out(430),
            product_re_out=>mul_re_out(430),
            product_im_out=>mul_im_out(430)
        );

    UMUL_431 : complex_multiplier
    generic map(
            re_multiplicator=>13538, --- 0.826293945312 + j-0.563171386719
            im_multiplicator=>-9227
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(431),
            data_im_in=>first_stage_im_out(431),
            product_re_out=>mul_re_out(431),
            product_im_out=>mul_im_out(431)
        );

    UMUL_432 : complex_multiplier
    generic map(
            re_multiplicator=>13159, --- 0.803161621094 + j-0.595642089844
            im_multiplicator=>-9759
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(432),
            data_im_in=>first_stage_im_out(432),
            product_re_out=>mul_re_out(432),
            product_im_out=>mul_im_out(432)
        );

    UMUL_433 : complex_multiplier
    generic map(
            re_multiplicator=>12760, --- 0.77880859375 + j-0.627197265625
            im_multiplicator=>-10276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(433),
            data_im_in=>first_stage_im_out(433),
            product_re_out=>mul_re_out(433),
            product_im_out=>mul_im_out(433)
        );

    UMUL_434 : complex_multiplier
    generic map(
            re_multiplicator=>12340, --- 0.753173828125 + j-0.657775878906
            im_multiplicator=>-10777
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(434),
            data_im_in=>first_stage_im_out(434),
            product_re_out=>mul_re_out(434),
            product_im_out=>mul_im_out(434)
        );

    UMUL_435 : complex_multiplier
    generic map(
            re_multiplicator=>11900, --- 0.726318359375 + j-0.687255859375
            im_multiplicator=>-11260
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(435),
            data_im_in=>first_stage_im_out(435),
            product_re_out=>mul_re_out(435),
            product_im_out=>mul_im_out(435)
        );

    UMUL_436 : complex_multiplier
    generic map(
            re_multiplicator=>11442, --- 0.698364257812 + j-0.715698242188
            im_multiplicator=>-11726
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(436),
            data_im_in=>first_stage_im_out(436),
            product_re_out=>mul_re_out(436),
            product_im_out=>mul_im_out(436)
        );

    UMUL_437 : complex_multiplier
    generic map(
            re_multiplicator=>10965, --- 0.669250488281 + j-0.742980957031
            im_multiplicator=>-12173
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(437),
            data_im_in=>first_stage_im_out(437),
            product_re_out=>mul_re_out(437),
            product_im_out=>mul_im_out(437)
        );

    UMUL_438 : complex_multiplier
    generic map(
            re_multiplicator=>10471, --- 0.639099121094 + j-0.76904296875
            im_multiplicator=>-12600
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(438),
            data_im_in=>first_stage_im_out(438),
            product_re_out=>mul_re_out(438),
            product_im_out=>mul_im_out(438)
        );

    UMUL_439 : complex_multiplier
    generic map(
            re_multiplicator=>9960, --- 0.60791015625 + j-0.7939453125
            im_multiplicator=>-13008
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(439),
            data_im_in=>first_stage_im_out(439),
            product_re_out=>mul_re_out(439),
            product_im_out=>mul_im_out(439)
        );

    UMUL_440 : complex_multiplier
    generic map(
            re_multiplicator=>9434, --- 0.575805664062 + j-0.817565917969
            im_multiplicator=>-13395
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(440),
            data_im_in=>first_stage_im_out(440),
            product_re_out=>mul_re_out(440),
            product_im_out=>mul_im_out(440)
        );

    UMUL_441 : complex_multiplier
    generic map(
            re_multiplicator=>8892, --- 0.542724609375 + j-0.83984375
            im_multiplicator=>-13760
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(441),
            data_im_in=>first_stage_im_out(441),
            product_re_out=>mul_re_out(441),
            product_im_out=>mul_im_out(441)
        );

    UMUL_442 : complex_multiplier
    generic map(
            re_multiplicator=>8336, --- 0.5087890625 + j-0.86083984375
            im_multiplicator=>-14104
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(442),
            data_im_in=>first_stage_im_out(442),
            product_re_out=>mul_re_out(442),
            product_im_out=>mul_im_out(442)
        );

    UMUL_443 : complex_multiplier
    generic map(
            re_multiplicator=>7767, --- 0.474060058594 + j-0.880432128906
            im_multiplicator=>-14425
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(443),
            data_im_in=>first_stage_im_out(443),
            product_re_out=>mul_re_out(443),
            product_im_out=>mul_im_out(443)
        );

    UMUL_444 : complex_multiplier
    generic map(
            re_multiplicator=>7186, --- 0.438598632812 + j-0.898620605469
            im_multiplicator=>-14723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(444),
            data_im_in=>first_stage_im_out(444),
            product_re_out=>mul_re_out(444),
            product_im_out=>mul_im_out(444)
        );

    UMUL_445 : complex_multiplier
    generic map(
            re_multiplicator=>6593, --- 0.402404785156 + j-0.915405273438
            im_multiplicator=>-14998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(445),
            data_im_in=>first_stage_im_out(445),
            product_re_out=>mul_re_out(445),
            product_im_out=>mul_im_out(445)
        );

    UMUL_446 : complex_multiplier
    generic map(
            re_multiplicator=>5990, --- 0.365600585938 + j-0.930725097656
            im_multiplicator=>-15249
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(446),
            data_im_in=>first_stage_im_out(446),
            product_re_out=>mul_re_out(446),
            product_im_out=>mul_im_out(446)
        );

    UMUL_447 : complex_multiplier
    generic map(
            re_multiplicator=>5377, --- 0.328186035156 + j-0.944580078125
            im_multiplicator=>-15476
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(447),
            data_im_in=>first_stage_im_out(447),
            product_re_out=>mul_re_out(447),
            product_im_out=>mul_im_out(447)
        );

    UDELAY_448_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(448),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(448)
        );
    UDELAY_448_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(448),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(448)
        );
    USHIFTER_448_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(448),
            data_out=>mul_re_out(448)
        );
    USHIFTER_448_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(448),
            data_out=>mul_im_out(448)
        );

    UMUL_449 : complex_multiplier
    generic map(
            re_multiplicator=>16368, --- 0.9990234375 + j-0.0429077148438
            im_multiplicator=>-703
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(449),
            data_im_in=>first_stage_im_out(449),
            product_re_out=>mul_re_out(449),
            product_im_out=>mul_im_out(449)
        );

    UMUL_450 : complex_multiplier
    generic map(
            re_multiplicator=>16323, --- 0.996276855469 + j-0.0857543945312
            im_multiplicator=>-1405
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(450),
            data_im_in=>first_stage_im_out(450),
            product_re_out=>mul_re_out(450),
            product_im_out=>mul_im_out(450)
        );

    UMUL_451 : complex_multiplier
    generic map(
            re_multiplicator=>16248, --- 0.99169921875 + j-0.128479003906
            im_multiplicator=>-2105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(451),
            data_im_in=>first_stage_im_out(451),
            product_re_out=>mul_re_out(451),
            product_im_out=>mul_im_out(451)
        );

    UMUL_452 : complex_multiplier
    generic map(
            re_multiplicator=>16142, --- 0.985229492188 + j-0.170959472656
            im_multiplicator=>-2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(452),
            data_im_in=>first_stage_im_out(452),
            product_re_out=>mul_re_out(452),
            product_im_out=>mul_im_out(452)
        );

    UMUL_453 : complex_multiplier
    generic map(
            re_multiplicator=>16007, --- 0.976989746094 + j-0.213073730469
            im_multiplicator=>-3491
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(453),
            data_im_in=>first_stage_im_out(453),
            product_re_out=>mul_re_out(453),
            product_im_out=>mul_im_out(453)
        );

    UMUL_454 : complex_multiplier
    generic map(
            re_multiplicator=>15842, --- 0.966918945312 + j-0.254821777344
            im_multiplicator=>-4175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(454),
            data_im_in=>first_stage_im_out(454),
            product_re_out=>mul_re_out(454),
            product_im_out=>mul_im_out(454)
        );

    UMUL_455 : complex_multiplier
    generic map(
            re_multiplicator=>15649, --- 0.955139160156 + j-0.296142578125
            im_multiplicator=>-4852
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(455),
            data_im_in=>first_stage_im_out(455),
            product_re_out=>mul_re_out(455),
            product_im_out=>mul_im_out(455)
        );

    UMUL_456 : complex_multiplier
    generic map(
            re_multiplicator=>15426, --- 0.941528320312 + j-0.336853027344
            im_multiplicator=>-5519
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(456),
            data_im_in=>first_stage_im_out(456),
            product_re_out=>mul_re_out(456),
            product_im_out=>mul_im_out(456)
        );

    UMUL_457 : complex_multiplier
    generic map(
            re_multiplicator=>15175, --- 0.926208496094 + j-0.376953125
            im_multiplicator=>-6176
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(457),
            data_im_in=>first_stage_im_out(457),
            product_re_out=>mul_re_out(457),
            product_im_out=>mul_im_out(457)
        );

    UMUL_458 : complex_multiplier
    generic map(
            re_multiplicator=>14895, --- 0.909118652344 + j-0.416381835938
            im_multiplicator=>-6822
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(458),
            data_im_in=>first_stage_im_out(458),
            product_re_out=>mul_re_out(458),
            product_im_out=>mul_im_out(458)
        );

    UMUL_459 : complex_multiplier
    generic map(
            re_multiplicator=>14589, --- 0.890441894531 + j-0.455078125
            im_multiplicator=>-7456
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(459),
            data_im_in=>first_stage_im_out(459),
            product_re_out=>mul_re_out(459),
            product_im_out=>mul_im_out(459)
        );

    UMUL_460 : complex_multiplier
    generic map(
            re_multiplicator=>14255, --- 0.870056152344 + j-0.492858886719
            im_multiplicator=>-8075
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(460),
            data_im_in=>first_stage_im_out(460),
            product_re_out=>mul_re_out(460),
            product_im_out=>mul_im_out(460)
        );

    UMUL_461 : complex_multiplier
    generic map(
            re_multiplicator=>13895, --- 0.848083496094 + j-0.52978515625
            im_multiplicator=>-8680
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(461),
            data_im_in=>first_stage_im_out(461),
            product_re_out=>mul_re_out(461),
            product_im_out=>mul_im_out(461)
        );

    UMUL_462 : complex_multiplier
    generic map(
            re_multiplicator=>13510, --- 0.824584960938 + j-0.565673828125
            im_multiplicator=>-9268
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(462),
            data_im_in=>first_stage_im_out(462),
            product_re_out=>mul_re_out(462),
            product_im_out=>mul_im_out(462)
        );

    UMUL_463 : complex_multiplier
    generic map(
            re_multiplicator=>13099, --- 0.799499511719 + j-0.6005859375
            im_multiplicator=>-9840
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(463),
            data_im_in=>first_stage_im_out(463),
            product_re_out=>mul_re_out(463),
            product_im_out=>mul_im_out(463)
        );

    UMUL_464 : complex_multiplier
    generic map(
            re_multiplicator=>12665, --- 0.773010253906 + j-0.634338378906
            im_multiplicator=>-10393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(464),
            data_im_in=>first_stage_im_out(464),
            product_re_out=>mul_re_out(464),
            product_im_out=>mul_im_out(464)
        );

    UMUL_465 : complex_multiplier
    generic map(
            re_multiplicator=>12207, --- 0.745056152344 + j-0.6669921875
            im_multiplicator=>-10928
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(465),
            data_im_in=>first_stage_im_out(465),
            product_re_out=>mul_re_out(465),
            product_im_out=>mul_im_out(465)
        );

    UMUL_466 : complex_multiplier
    generic map(
            re_multiplicator=>11726, --- 0.715698242188 + j-0.698364257812
            im_multiplicator=>-11442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(466),
            data_im_in=>first_stage_im_out(466),
            product_re_out=>mul_re_out(466),
            product_im_out=>mul_im_out(466)
        );

    UMUL_467 : complex_multiplier
    generic map(
            re_multiplicator=>11224, --- 0.68505859375 + j-0.728454589844
            im_multiplicator=>-11935
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(467),
            data_im_in=>first_stage_im_out(467),
            product_re_out=>mul_re_out(467),
            product_im_out=>mul_im_out(467)
        );

    UMUL_468 : complex_multiplier
    generic map(
            re_multiplicator=>10701, --- 0.653137207031 + j-0.757202148438
            im_multiplicator=>-12406
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(468),
            data_im_in=>first_stage_im_out(468),
            product_re_out=>mul_re_out(468),
            product_im_out=>mul_im_out(468)
        );

    UMUL_469 : complex_multiplier
    generic map(
            re_multiplicator=>10159, --- 0.620056152344 + j-0.784545898438
            im_multiplicator=>-12854
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(469),
            data_im_in=>first_stage_im_out(469),
            product_re_out=>mul_re_out(469),
            product_im_out=>mul_im_out(469)
        );

    UMUL_470 : complex_multiplier
    generic map(
            re_multiplicator=>9597, --- 0.585754394531 + j-0.810424804688
            im_multiplicator=>-13278
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(470),
            data_im_in=>first_stage_im_out(470),
            product_re_out=>mul_re_out(470),
            product_im_out=>mul_im_out(470)
        );

    UMUL_471 : complex_multiplier
    generic map(
            re_multiplicator=>9018, --- 0.550415039062 + j-0.834838867188
            im_multiplicator=>-13678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(471),
            data_im_in=>first_stage_im_out(471),
            product_re_out=>mul_re_out(471),
            product_im_out=>mul_im_out(471)
        );

    UMUL_472 : complex_multiplier
    generic map(
            re_multiplicator=>8423, --- 0.514099121094 + j-0.857727050781
            im_multiplicator=>-14053
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(472),
            data_im_in=>first_stage_im_out(472),
            product_re_out=>mul_re_out(472),
            product_im_out=>mul_im_out(472)
        );

    UMUL_473 : complex_multiplier
    generic map(
            re_multiplicator=>7811, --- 0.476745605469 + j-0.878967285156
            im_multiplicator=>-14401
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(473),
            data_im_in=>first_stage_im_out(473),
            product_re_out=>mul_re_out(473),
            product_im_out=>mul_im_out(473)
        );

    UMUL_474 : complex_multiplier
    generic map(
            re_multiplicator=>7186, --- 0.438598632812 + j-0.898620605469
            im_multiplicator=>-14723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(474),
            data_im_in=>first_stage_im_out(474),
            product_re_out=>mul_re_out(474),
            product_im_out=>mul_im_out(474)
        );

    UMUL_475 : complex_multiplier
    generic map(
            re_multiplicator=>6547, --- 0.399597167969 + j-0.916625976562
            im_multiplicator=>-15018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(475),
            data_im_in=>first_stage_im_out(475),
            product_re_out=>mul_re_out(475),
            product_im_out=>mul_im_out(475)
        );

    UMUL_476 : complex_multiplier
    generic map(
            re_multiplicator=>5896, --- 0.35986328125 + j-0.932983398438
            im_multiplicator=>-15286
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(476),
            data_im_in=>first_stage_im_out(476),
            product_re_out=>mul_re_out(476),
            product_im_out=>mul_im_out(476)
        );

    UMUL_477 : complex_multiplier
    generic map(
            re_multiplicator=>5234, --- 0.319458007812 + j-0.947570800781
            im_multiplicator=>-15525
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(477),
            data_im_in=>first_stage_im_out(477),
            product_re_out=>mul_re_out(477),
            product_im_out=>mul_im_out(477)
        );

    UMUL_478 : complex_multiplier
    generic map(
            re_multiplicator=>4563, --- 0.278503417969 + j-0.960388183594
            im_multiplicator=>-15735
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(478),
            data_im_in=>first_stage_im_out(478),
            product_re_out=>mul_re_out(478),
            product_im_out=>mul_im_out(478)
        );

    UMUL_479 : complex_multiplier
    generic map(
            re_multiplicator=>3883, --- 0.236999511719 + j-0.971496582031
            im_multiplicator=>-15917
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(479),
            data_im_in=>first_stage_im_out(479),
            product_re_out=>mul_re_out(479),
            product_im_out=>mul_im_out(479)
        );

    UDELAY_480_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(480),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(480)
        );
    UDELAY_480_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(480),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(480)
        );
    USHIFTER_480_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(480),
            data_out=>mul_re_out(480)
        );
    USHIFTER_480_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(480),
            data_out=>mul_im_out(480)
        );

    UMUL_481 : complex_multiplier
    generic map(
            re_multiplicator=>16366, --- 0.998901367188 + j-0.0459594726562
            im_multiplicator=>-753
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(481),
            data_im_in=>first_stage_im_out(481),
            product_re_out=>mul_re_out(481),
            product_im_out=>mul_im_out(481)
        );

    UMUL_482 : complex_multiplier
    generic map(
            re_multiplicator=>16314, --- 0.995727539062 + j-0.0918579101562
            im_multiplicator=>-1505
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(482),
            data_im_in=>first_stage_im_out(482),
            product_re_out=>mul_re_out(482),
            product_im_out=>mul_im_out(482)
        );

    UMUL_483 : complex_multiplier
    generic map(
            re_multiplicator=>16228, --- 0.990478515625 + j-0.137573242188
            im_multiplicator=>-2254
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(483),
            data_im_in=>first_stage_im_out(483),
            product_re_out=>mul_re_out(483),
            product_im_out=>mul_im_out(483)
        );

    UMUL_484 : complex_multiplier
    generic map(
            re_multiplicator=>16107, --- 0.983093261719 + j-0.182983398438
            im_multiplicator=>-2998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(484),
            data_im_in=>first_stage_im_out(484),
            product_re_out=>mul_re_out(484),
            product_im_out=>mul_im_out(484)
        );

    UMUL_485 : complex_multiplier
    generic map(
            re_multiplicator=>15952, --- 0.9736328125 + j-0.22802734375
            im_multiplicator=>-3736
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(485),
            data_im_in=>first_stage_im_out(485),
            product_re_out=>mul_re_out(485),
            product_im_out=>mul_im_out(485)
        );

    UMUL_486 : complex_multiplier
    generic map(
            re_multiplicator=>15763, --- 0.962097167969 + j-0.272583007812
            im_multiplicator=>-4466
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(486),
            data_im_in=>first_stage_im_out(486),
            product_re_out=>mul_re_out(486),
            product_im_out=>mul_im_out(486)
        );

    UMUL_487 : complex_multiplier
    generic map(
            re_multiplicator=>15541, --- 0.948547363281 + j-0.316589355469
            im_multiplicator=>-5187
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(487),
            data_im_in=>first_stage_im_out(487),
            product_re_out=>mul_re_out(487),
            product_im_out=>mul_im_out(487)
        );

    UMUL_488 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(488),
            data_im_in=>first_stage_im_out(488),
            product_re_out=>mul_re_out(488),
            product_im_out=>mul_im_out(488)
        );

    UMUL_489 : complex_multiplier
    generic map(
            re_multiplicator=>14998, --- 0.915405273438 + j-0.402404785156
            im_multiplicator=>-6593
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(489),
            data_im_in=>first_stage_im_out(489),
            product_re_out=>mul_re_out(489),
            product_im_out=>mul_im_out(489)
        );

    UMUL_490 : complex_multiplier
    generic map(
            re_multiplicator=>14679, --- 0.895935058594 + j-0.444091796875
            im_multiplicator=>-7276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(490),
            data_im_in=>first_stage_im_out(490),
            product_re_out=>mul_re_out(490),
            product_im_out=>mul_im_out(490)
        );

    UMUL_491 : complex_multiplier
    generic map(
            re_multiplicator=>14329, --- 0.874572753906 + j-0.48486328125
            im_multiplicator=>-7944
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(491),
            data_im_in=>first_stage_im_out(491),
            product_re_out=>mul_re_out(491),
            product_im_out=>mul_im_out(491)
        );

    UMUL_492 : complex_multiplier
    generic map(
            re_multiplicator=>13948, --- 0.851318359375 + j-0.524536132812
            im_multiplicator=>-8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(492),
            data_im_in=>first_stage_im_out(492),
            product_re_out=>mul_re_out(492),
            product_im_out=>mul_im_out(492)
        );

    UMUL_493 : complex_multiplier
    generic map(
            re_multiplicator=>13538, --- 0.826293945312 + j-0.563171386719
            im_multiplicator=>-9227
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(493),
            data_im_in=>first_stage_im_out(493),
            product_re_out=>mul_re_out(493),
            product_im_out=>mul_im_out(493)
        );

    UMUL_494 : complex_multiplier
    generic map(
            re_multiplicator=>13099, --- 0.799499511719 + j-0.6005859375
            im_multiplicator=>-9840
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(494),
            data_im_in=>first_stage_im_out(494),
            product_re_out=>mul_re_out(494),
            product_im_out=>mul_im_out(494)
        );

    UMUL_495 : complex_multiplier
    generic map(
            re_multiplicator=>12633, --- 0.771057128906 + j-0.63671875
            im_multiplicator=>-10432
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(495),
            data_im_in=>first_stage_im_out(495),
            product_re_out=>mul_re_out(495),
            product_im_out=>mul_im_out(495)
        );

    UMUL_496 : complex_multiplier
    generic map(
            re_multiplicator=>12139, --- 0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(496),
            data_im_in=>first_stage_im_out(496),
            product_re_out=>mul_re_out(496),
            product_im_out=>mul_im_out(496)
        );

    UMUL_497 : complex_multiplier
    generic map(
            re_multiplicator=>11620, --- 0.709228515625 + j-0.704895019531
            im_multiplicator=>-11549
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(497),
            data_im_in=>first_stage_im_out(497),
            product_re_out=>mul_re_out(497),
            product_im_out=>mul_im_out(497)
        );

    UMUL_498 : complex_multiplier
    generic map(
            re_multiplicator=>11077, --- 0.676086425781 + j-0.73681640625
            im_multiplicator=>-12072
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(498),
            data_im_in=>first_stage_im_out(498),
            product_re_out=>mul_re_out(498),
            product_im_out=>mul_im_out(498)
        );

    UMUL_499 : complex_multiplier
    generic map(
            re_multiplicator=>10510, --- 0.641479492188 + j-0.76708984375
            im_multiplicator=>-12568
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(499),
            data_im_in=>first_stage_im_out(499),
            product_re_out=>mul_re_out(499),
            product_im_out=>mul_im_out(499)
        );

    UMUL_500 : complex_multiplier
    generic map(
            re_multiplicator=>9920, --- 0.60546875 + j-0.795776367188
            im_multiplicator=>-13038
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(500),
            data_im_in=>first_stage_im_out(500),
            product_re_out=>mul_re_out(500),
            product_im_out=>mul_im_out(500)
        );

    UMUL_501 : complex_multiplier
    generic map(
            re_multiplicator=>9310, --- 0.568237304688 + j-0.822814941406
            im_multiplicator=>-13481
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(501),
            data_im_in=>first_stage_im_out(501),
            product_re_out=>mul_re_out(501),
            product_im_out=>mul_im_out(501)
        );

    UMUL_502 : complex_multiplier
    generic map(
            re_multiplicator=>8680, --- 0.52978515625 + j-0.848083496094
            im_multiplicator=>-13895
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(502),
            data_im_in=>first_stage_im_out(502),
            product_re_out=>mul_re_out(502),
            product_im_out=>mul_im_out(502)
        );

    UMUL_503 : complex_multiplier
    generic map(
            re_multiplicator=>8031, --- 0.490173339844 + j-0.87158203125
            im_multiplicator=>-14280
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(503),
            data_im_in=>first_stage_im_out(503),
            product_re_out=>mul_re_out(503),
            product_im_out=>mul_im_out(503)
        );

    UMUL_504 : complex_multiplier
    generic map(
            re_multiplicator=>7366, --- 0.449584960938 + j-0.893188476562
            im_multiplicator=>-14634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(504),
            data_im_in=>first_stage_im_out(504),
            product_re_out=>mul_re_out(504),
            product_im_out=>mul_im_out(504)
        );

    UMUL_505 : complex_multiplier
    generic map(
            re_multiplicator=>6685, --- 0.408020019531 + j-0.912902832031
            im_multiplicator=>-14957
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(505),
            data_im_in=>first_stage_im_out(505),
            product_re_out=>mul_re_out(505),
            product_im_out=>mul_im_out(505)
        );

    UMUL_506 : complex_multiplier
    generic map(
            re_multiplicator=>5990, --- 0.365600585938 + j-0.930725097656
            im_multiplicator=>-15249
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(506),
            data_im_in=>first_stage_im_out(506),
            product_re_out=>mul_re_out(506),
            product_im_out=>mul_im_out(506)
        );

    UMUL_507 : complex_multiplier
    generic map(
            re_multiplicator=>5282, --- 0.322387695312 + j-0.946594238281
            im_multiplicator=>-15509
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(507),
            data_im_in=>first_stage_im_out(507),
            product_re_out=>mul_re_out(507),
            product_im_out=>mul_im_out(507)
        );

    UMUL_508 : complex_multiplier
    generic map(
            re_multiplicator=>4563, --- 0.278503417969 + j-0.960388183594
            im_multiplicator=>-15735
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(508),
            data_im_in=>first_stage_im_out(508),
            product_re_out=>mul_re_out(508),
            product_im_out=>mul_im_out(508)
        );

    UMUL_509 : complex_multiplier
    generic map(
            re_multiplicator=>3834, --- 0.234008789062 + j-0.97216796875
            im_multiplicator=>-15928
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(509),
            data_im_in=>first_stage_im_out(509),
            product_re_out=>mul_re_out(509),
            product_im_out=>mul_im_out(509)
        );

    UMUL_510 : complex_multiplier
    generic map(
            re_multiplicator=>3097, --- 0.189025878906 + j-0.98193359375
            im_multiplicator=>-16088
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(510),
            data_im_in=>first_stage_im_out(510),
            product_re_out=>mul_re_out(510),
            product_im_out=>mul_im_out(510)
        );

    UMUL_511 : complex_multiplier
    generic map(
            re_multiplicator=>2354, --- 0.143676757812 + j-0.989562988281
            im_multiplicator=>-16213
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(511),
            data_im_in=>first_stage_im_out(511),
            product_re_out=>mul_re_out(511),
            product_im_out=>mul_im_out(511)
        );

    UDELAY_512_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(512),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(512)
        );
    UDELAY_512_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(512),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(512)
        );
    USHIFTER_512_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(512),
            data_out=>mul_re_out(512)
        );
    USHIFTER_512_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(512),
            data_out=>mul_im_out(512)
        );

    UMUL_513 : complex_multiplier
    generic map(
            re_multiplicator=>16364, --- 0.998779296875 + j-0.0490112304688
            im_multiplicator=>-803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(513),
            data_im_in=>first_stage_im_out(513),
            product_re_out=>mul_re_out(513),
            product_im_out=>mul_im_out(513)
        );

    UMUL_514 : complex_multiplier
    generic map(
            re_multiplicator=>16305, --- 0.995178222656 + j-0.0979614257812
            im_multiplicator=>-1605
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(514),
            data_im_in=>first_stage_im_out(514),
            product_re_out=>mul_re_out(514),
            product_im_out=>mul_im_out(514)
        );

    UMUL_515 : complex_multiplier
    generic map(
            re_multiplicator=>16206, --- 0.989135742188 + j-0.146728515625
            im_multiplicator=>-2404
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(515),
            data_im_in=>first_stage_im_out(515),
            product_re_out=>mul_re_out(515),
            product_im_out=>mul_im_out(515)
        );

    UMUL_516 : complex_multiplier
    generic map(
            re_multiplicator=>16069, --- 0.980773925781 + j-0.195068359375
            im_multiplicator=>-3196
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(516),
            data_im_in=>first_stage_im_out(516),
            product_re_out=>mul_re_out(516),
            product_im_out=>mul_im_out(516)
        );

    UMUL_517 : complex_multiplier
    generic map(
            re_multiplicator=>15892, --- 0.969970703125 + j-0.242919921875
            im_multiplicator=>-3980
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(517),
            data_im_in=>first_stage_im_out(517),
            product_re_out=>mul_re_out(517),
            product_im_out=>mul_im_out(517)
        );

    UMUL_518 : complex_multiplier
    generic map(
            re_multiplicator=>15678, --- 0.956909179688 + j-0.290283203125
            im_multiplicator=>-4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(518),
            data_im_in=>first_stage_im_out(518),
            product_re_out=>mul_re_out(518),
            product_im_out=>mul_im_out(518)
        );

    UMUL_519 : complex_multiplier
    generic map(
            re_multiplicator=>15426, --- 0.941528320312 + j-0.336853027344
            im_multiplicator=>-5519
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(519),
            data_im_in=>first_stage_im_out(519),
            product_re_out=>mul_re_out(519),
            product_im_out=>mul_im_out(519)
        );

    UMUL_520 : complex_multiplier
    generic map(
            re_multiplicator=>15136, --- 0.923828125 + j-0.382629394531
            im_multiplicator=>-6269
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(520),
            data_im_in=>first_stage_im_out(520),
            product_re_out=>mul_re_out(520),
            product_im_out=>mul_im_out(520)
        );

    UMUL_521 : complex_multiplier
    generic map(
            re_multiplicator=>14810, --- 0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(521),
            data_im_in=>first_stage_im_out(521),
            product_re_out=>mul_re_out(521),
            product_im_out=>mul_im_out(521)
        );

    UMUL_522 : complex_multiplier
    generic map(
            re_multiplicator=>14449, --- 0.881896972656 + j-0.471374511719
            im_multiplicator=>-7723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(522),
            data_im_in=>first_stage_im_out(522),
            product_re_out=>mul_re_out(522),
            product_im_out=>mul_im_out(522)
        );

    UMUL_523 : complex_multiplier
    generic map(
            re_multiplicator=>14053, --- 0.857727050781 + j-0.514099121094
            im_multiplicator=>-8423
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(523),
            data_im_in=>first_stage_im_out(523),
            product_re_out=>mul_re_out(523),
            product_im_out=>mul_im_out(523)
        );

    UMUL_524 : complex_multiplier
    generic map(
            re_multiplicator=>13622, --- 0.831420898438 + j-0.555541992188
            im_multiplicator=>-9102
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(524),
            data_im_in=>first_stage_im_out(524),
            product_re_out=>mul_re_out(524),
            product_im_out=>mul_im_out(524)
        );

    UMUL_525 : complex_multiplier
    generic map(
            re_multiplicator=>13159, --- 0.803161621094 + j-0.595642089844
            im_multiplicator=>-9759
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(525),
            data_im_in=>first_stage_im_out(525),
            product_re_out=>mul_re_out(525),
            product_im_out=>mul_im_out(525)
        );

    UMUL_526 : complex_multiplier
    generic map(
            re_multiplicator=>12665, --- 0.773010253906 + j-0.634338378906
            im_multiplicator=>-10393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(526),
            data_im_in=>first_stage_im_out(526),
            product_re_out=>mul_re_out(526),
            product_im_out=>mul_im_out(526)
        );

    UMUL_527 : complex_multiplier
    generic map(
            re_multiplicator=>12139, --- 0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(527),
            data_im_in=>first_stage_im_out(527),
            product_re_out=>mul_re_out(527),
            product_im_out=>mul_im_out(527)
        );

    UMUL_528 : complex_multiplier
    generic map(
            re_multiplicator=>11585, --- 0.707092285156 + j-0.707092285156
            im_multiplicator=>-11585
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(528),
            data_im_in=>first_stage_im_out(528),
            product_re_out=>mul_re_out(528),
            product_im_out=>mul_im_out(528)
        );

    UMUL_529 : complex_multiplier
    generic map(
            re_multiplicator=>11002, --- 0.671508789062 + j-0.740905761719
            im_multiplicator=>-12139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(529),
            data_im_in=>first_stage_im_out(529),
            product_re_out=>mul_re_out(529),
            product_im_out=>mul_im_out(529)
        );

    UMUL_530 : complex_multiplier
    generic map(
            re_multiplicator=>10393, --- 0.634338378906 + j-0.773010253906
            im_multiplicator=>-12665
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(530),
            data_im_in=>first_stage_im_out(530),
            product_re_out=>mul_re_out(530),
            product_im_out=>mul_im_out(530)
        );

    UMUL_531 : complex_multiplier
    generic map(
            re_multiplicator=>9759, --- 0.595642089844 + j-0.803161621094
            im_multiplicator=>-13159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(531),
            data_im_in=>first_stage_im_out(531),
            product_re_out=>mul_re_out(531),
            product_im_out=>mul_im_out(531)
        );

    UMUL_532 : complex_multiplier
    generic map(
            re_multiplicator=>9102, --- 0.555541992188 + j-0.831420898438
            im_multiplicator=>-13622
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(532),
            data_im_in=>first_stage_im_out(532),
            product_re_out=>mul_re_out(532),
            product_im_out=>mul_im_out(532)
        );

    UMUL_533 : complex_multiplier
    generic map(
            re_multiplicator=>8423, --- 0.514099121094 + j-0.857727050781
            im_multiplicator=>-14053
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(533),
            data_im_in=>first_stage_im_out(533),
            product_re_out=>mul_re_out(533),
            product_im_out=>mul_im_out(533)
        );

    UMUL_534 : complex_multiplier
    generic map(
            re_multiplicator=>7723, --- 0.471374511719 + j-0.881896972656
            im_multiplicator=>-14449
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(534),
            data_im_in=>first_stage_im_out(534),
            product_re_out=>mul_re_out(534),
            product_im_out=>mul_im_out(534)
        );

    UMUL_535 : complex_multiplier
    generic map(
            re_multiplicator=>7005, --- 0.427551269531 + j-0.903930664062
            im_multiplicator=>-14810
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(535),
            data_im_in=>first_stage_im_out(535),
            product_re_out=>mul_re_out(535),
            product_im_out=>mul_im_out(535)
        );

    UMUL_536 : complex_multiplier
    generic map(
            re_multiplicator=>6269, --- 0.382629394531 + j-0.923828125
            im_multiplicator=>-15136
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(536),
            data_im_in=>first_stage_im_out(536),
            product_re_out=>mul_re_out(536),
            product_im_out=>mul_im_out(536)
        );

    UMUL_537 : complex_multiplier
    generic map(
            re_multiplicator=>5519, --- 0.336853027344 + j-0.941528320312
            im_multiplicator=>-15426
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(537),
            data_im_in=>first_stage_im_out(537),
            product_re_out=>mul_re_out(537),
            product_im_out=>mul_im_out(537)
        );

    UMUL_538 : complex_multiplier
    generic map(
            re_multiplicator=>4756, --- 0.290283203125 + j-0.956909179688
            im_multiplicator=>-15678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(538),
            data_im_in=>first_stage_im_out(538),
            product_re_out=>mul_re_out(538),
            product_im_out=>mul_im_out(538)
        );

    UMUL_539 : complex_multiplier
    generic map(
            re_multiplicator=>3980, --- 0.242919921875 + j-0.969970703125
            im_multiplicator=>-15892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(539),
            data_im_in=>first_stage_im_out(539),
            product_re_out=>mul_re_out(539),
            product_im_out=>mul_im_out(539)
        );

    UMUL_540 : complex_multiplier
    generic map(
            re_multiplicator=>3196, --- 0.195068359375 + j-0.980773925781
            im_multiplicator=>-16069
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(540),
            data_im_in=>first_stage_im_out(540),
            product_re_out=>mul_re_out(540),
            product_im_out=>mul_im_out(540)
        );

    UMUL_541 : complex_multiplier
    generic map(
            re_multiplicator=>2404, --- 0.146728515625 + j-0.989135742188
            im_multiplicator=>-16206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(541),
            data_im_in=>first_stage_im_out(541),
            product_re_out=>mul_re_out(541),
            product_im_out=>mul_im_out(541)
        );

    UMUL_542 : complex_multiplier
    generic map(
            re_multiplicator=>1605, --- 0.0979614257812 + j-0.995178222656
            im_multiplicator=>-16305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(542),
            data_im_in=>first_stage_im_out(542),
            product_re_out=>mul_re_out(542),
            product_im_out=>mul_im_out(542)
        );

    UMUL_543 : complex_multiplier
    generic map(
            re_multiplicator=>803, --- 0.0490112304688 + j-0.998779296875
            im_multiplicator=>-16364
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(543),
            data_im_in=>first_stage_im_out(543),
            product_re_out=>mul_re_out(543),
            product_im_out=>mul_im_out(543)
        );

    UDELAY_544_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(544),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(544)
        );
    UDELAY_544_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(544),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(544)
        );
    USHIFTER_544_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(544),
            data_out=>mul_re_out(544)
        );
    USHIFTER_544_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(544),
            data_out=>mul_im_out(544)
        );

    UMUL_545 : complex_multiplier
    generic map(
            re_multiplicator=>16361, --- 0.998596191406 + j-0.0521240234375
            im_multiplicator=>-854
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(545),
            data_im_in=>first_stage_im_out(545),
            product_re_out=>mul_re_out(545),
            product_im_out=>mul_im_out(545)
        );

    UMUL_546 : complex_multiplier
    generic map(
            re_multiplicator=>16294, --- 0.994506835938 + j-0.104064941406
            im_multiplicator=>-1705
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(546),
            data_im_in=>first_stage_im_out(546),
            product_re_out=>mul_re_out(546),
            product_im_out=>mul_im_out(546)
        );

    UMUL_547 : complex_multiplier
    generic map(
            re_multiplicator=>16183, --- 0.987731933594 + j-0.155822753906
            im_multiplicator=>-2553
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(547),
            data_im_in=>first_stage_im_out(547),
            product_re_out=>mul_re_out(547),
            product_im_out=>mul_im_out(547)
        );

    UMUL_548 : complex_multiplier
    generic map(
            re_multiplicator=>16028, --- 0.978271484375 + j-0.207092285156
            im_multiplicator=>-3393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(548),
            data_im_in=>first_stage_im_out(548),
            product_re_out=>mul_re_out(548),
            product_im_out=>mul_im_out(548)
        );

    UMUL_549 : complex_multiplier
    generic map(
            re_multiplicator=>15830, --- 0.966186523438 + j-0.2578125
            im_multiplicator=>-4224
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(549),
            data_im_in=>first_stage_im_out(549),
            product_re_out=>mul_re_out(549),
            product_im_out=>mul_im_out(549)
        );

    UMUL_550 : complex_multiplier
    generic map(
            re_multiplicator=>15588, --- 0.951416015625 + j-0.307800292969
            im_multiplicator=>-5043
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(550),
            data_im_in=>first_stage_im_out(550),
            product_re_out=>mul_re_out(550),
            product_im_out=>mul_im_out(550)
        );

    UMUL_551 : complex_multiplier
    generic map(
            re_multiplicator=>15304, --- 0.93408203125 + j-0.356994628906
            im_multiplicator=>-5849
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(551),
            data_im_in=>first_stage_im_out(551),
            product_re_out=>mul_re_out(551),
            product_im_out=>mul_im_out(551)
        );

    UMUL_552 : complex_multiplier
    generic map(
            re_multiplicator=>14978, --- 0.914184570312 + j-0.405212402344
            im_multiplicator=>-6639
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(552),
            data_im_in=>first_stage_im_out(552),
            product_re_out=>mul_re_out(552),
            product_im_out=>mul_im_out(552)
        );

    UMUL_553 : complex_multiplier
    generic map(
            re_multiplicator=>14611, --- 0.891784667969 + j-0.452331542969
            im_multiplicator=>-7411
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(553),
            data_im_in=>first_stage_im_out(553),
            product_re_out=>mul_re_out(553),
            product_im_out=>mul_im_out(553)
        );

    UMUL_554 : complex_multiplier
    generic map(
            re_multiplicator=>14205, --- 0.867004394531 + j-0.498168945312
            im_multiplicator=>-8162
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(554),
            data_im_in=>first_stage_im_out(554),
            product_re_out=>mul_re_out(554),
            product_im_out=>mul_im_out(554)
        );

    UMUL_555 : complex_multiplier
    generic map(
            re_multiplicator=>13760, --- 0.83984375 + j-0.542724609375
            im_multiplicator=>-8892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(555),
            data_im_in=>first_stage_im_out(555),
            product_re_out=>mul_re_out(555),
            product_im_out=>mul_im_out(555)
        );

    UMUL_556 : complex_multiplier
    generic map(
            re_multiplicator=>13278, --- 0.810424804688 + j-0.585754394531
            im_multiplicator=>-9597
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(556),
            data_im_in=>first_stage_im_out(556),
            product_re_out=>mul_re_out(556),
            product_im_out=>mul_im_out(556)
        );

    UMUL_557 : complex_multiplier
    generic map(
            re_multiplicator=>12760, --- 0.77880859375 + j-0.627197265625
            im_multiplicator=>-10276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(557),
            data_im_in=>first_stage_im_out(557),
            product_re_out=>mul_re_out(557),
            product_im_out=>mul_im_out(557)
        );

    UMUL_558 : complex_multiplier
    generic map(
            re_multiplicator=>12207, --- 0.745056152344 + j-0.6669921875
            im_multiplicator=>-10928
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(558),
            data_im_in=>first_stage_im_out(558),
            product_re_out=>mul_re_out(558),
            product_im_out=>mul_im_out(558)
        );

    UMUL_559 : complex_multiplier
    generic map(
            re_multiplicator=>11620, --- 0.709228515625 + j-0.704895019531
            im_multiplicator=>-11549
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(559),
            data_im_in=>first_stage_im_out(559),
            product_re_out=>mul_re_out(559),
            product_im_out=>mul_im_out(559)
        );

    UMUL_560 : complex_multiplier
    generic map(
            re_multiplicator=>11002, --- 0.671508789062 + j-0.740905761719
            im_multiplicator=>-12139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(560),
            data_im_in=>first_stage_im_out(560),
            product_re_out=>mul_re_out(560),
            product_im_out=>mul_im_out(560)
        );

    UMUL_561 : complex_multiplier
    generic map(
            re_multiplicator=>10354, --- 0.631958007812 + j-0.77490234375
            im_multiplicator=>-12696
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(561),
            data_im_in=>first_stage_im_out(561),
            product_re_out=>mul_re_out(561),
            product_im_out=>mul_im_out(561)
        );

    UMUL_562 : complex_multiplier
    generic map(
            re_multiplicator=>9679, --- 0.590759277344 + j-0.806823730469
            im_multiplicator=>-13219
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(562),
            data_im_in=>first_stage_im_out(562),
            product_re_out=>mul_re_out(562),
            product_im_out=>mul_im_out(562)
        );

    UMUL_563 : complex_multiplier
    generic map(
            re_multiplicator=>8976, --- 0.5478515625 + j-0.836486816406
            im_multiplicator=>-13705
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(563),
            data_im_in=>first_stage_im_out(563),
            product_re_out=>mul_re_out(563),
            product_im_out=>mul_im_out(563)
        );

    UMUL_564 : complex_multiplier
    generic map(
            re_multiplicator=>8249, --- 0.503479003906 + j-0.863952636719
            im_multiplicator=>-14155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(564),
            data_im_in=>first_stage_im_out(564),
            product_re_out=>mul_re_out(564),
            product_im_out=>mul_im_out(564)
        );

    UMUL_565 : complex_multiplier
    generic map(
            re_multiplicator=>7500, --- 0.457763671875 + j-0.889038085938
            im_multiplicator=>-14566
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(565),
            data_im_in=>first_stage_im_out(565),
            product_re_out=>mul_re_out(565),
            product_im_out=>mul_im_out(565)
        );

    UMUL_566 : complex_multiplier
    generic map(
            re_multiplicator=>6731, --- 0.410827636719 + j-0.911682128906
            im_multiplicator=>-14937
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(566),
            data_im_in=>first_stage_im_out(566),
            product_re_out=>mul_re_out(566),
            product_im_out=>mul_im_out(566)
        );

    UMUL_567 : complex_multiplier
    generic map(
            re_multiplicator=>5943, --- 0.362731933594 + j-0.931823730469
            im_multiplicator=>-15267
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(567),
            data_im_in=>first_stage_im_out(567),
            product_re_out=>mul_re_out(567),
            product_im_out=>mul_im_out(567)
        );

    UMUL_568 : complex_multiplier
    generic map(
            re_multiplicator=>5139, --- 0.313659667969 + j-0.949523925781
            im_multiplicator=>-15557
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(568),
            data_im_in=>first_stage_im_out(568),
            product_re_out=>mul_re_out(568),
            product_im_out=>mul_im_out(568)
        );

    UMUL_569 : complex_multiplier
    generic map(
            re_multiplicator=>4321, --- 0.263732910156 + j-0.964538574219
            im_multiplicator=>-15803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(569),
            data_im_in=>first_stage_im_out(569),
            product_re_out=>mul_re_out(569),
            product_im_out=>mul_im_out(569)
        );

    UMUL_570 : complex_multiplier
    generic map(
            re_multiplicator=>3491, --- 0.213073730469 + j-0.976989746094
            im_multiplicator=>-16007
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(570),
            data_im_in=>first_stage_im_out(570),
            product_re_out=>mul_re_out(570),
            product_im_out=>mul_im_out(570)
        );

    UMUL_571 : complex_multiplier
    generic map(
            re_multiplicator=>2652, --- 0.161865234375 + j-0.986755371094
            im_multiplicator=>-16167
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(571),
            data_im_in=>first_stage_im_out(571),
            product_re_out=>mul_re_out(571),
            product_im_out=>mul_im_out(571)
        );

    UMUL_572 : complex_multiplier
    generic map(
            re_multiplicator=>1805, --- 0.110168457031 + j-0.993896484375
            im_multiplicator=>-16284
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(572),
            data_im_in=>first_stage_im_out(572),
            product_re_out=>mul_re_out(572),
            product_im_out=>mul_im_out(572)
        );

    UMUL_573 : complex_multiplier
    generic map(
            re_multiplicator=>954, --- 0.0582275390625 + j-0.998291015625
            im_multiplicator=>-16356
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(573),
            data_im_in=>first_stage_im_out(573),
            product_re_out=>mul_re_out(573),
            product_im_out=>mul_im_out(573)
        );

    UMUL_574 : complex_multiplier
    generic map(
            re_multiplicator=>100, --- 0.006103515625 + j-0.999938964844
            im_multiplicator=>-16383
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(574),
            data_im_in=>first_stage_im_out(574),
            product_re_out=>mul_re_out(574),
            product_im_out=>mul_im_out(574)
        );

    UMUL_575 : complex_multiplier
    generic map(
            re_multiplicator=>-753, --- -0.0459594726562 + j-0.998901367188
            im_multiplicator=>-16366
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(575),
            data_im_in=>first_stage_im_out(575),
            product_re_out=>mul_re_out(575),
            product_im_out=>mul_im_out(575)
        );

    UDELAY_576_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(576),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(576)
        );
    UDELAY_576_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(576),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(576)
        );
    USHIFTER_576_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(576),
            data_out=>mul_re_out(576)
        );
    USHIFTER_576_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(576),
            data_out=>mul_im_out(576)
        );

    UMUL_577 : complex_multiplier
    generic map(
            re_multiplicator=>16359, --- 0.998474121094 + j-0.05517578125
            im_multiplicator=>-904
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(577),
            data_im_in=>first_stage_im_out(577),
            product_re_out=>mul_re_out(577),
            product_im_out=>mul_im_out(577)
        );

    UMUL_578 : complex_multiplier
    generic map(
            re_multiplicator=>16284, --- 0.993896484375 + j-0.110168457031
            im_multiplicator=>-1805
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(578),
            data_im_in=>first_stage_im_out(578),
            product_re_out=>mul_re_out(578),
            product_im_out=>mul_im_out(578)
        );

    UMUL_579 : complex_multiplier
    generic map(
            re_multiplicator=>16159, --- 0.986267089844 + j-0.164855957031
            im_multiplicator=>-2701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(579),
            data_im_in=>first_stage_im_out(579),
            product_re_out=>mul_re_out(579),
            product_im_out=>mul_im_out(579)
        );

    UMUL_580 : complex_multiplier
    generic map(
            re_multiplicator=>15985, --- 0.975646972656 + j-0.219055175781
            im_multiplicator=>-3589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(580),
            data_im_in=>first_stage_im_out(580),
            product_re_out=>mul_re_out(580),
            product_im_out=>mul_im_out(580)
        );

    UMUL_581 : complex_multiplier
    generic map(
            re_multiplicator=>15763, --- 0.962097167969 + j-0.272583007812
            im_multiplicator=>-4466
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(581),
            data_im_in=>first_stage_im_out(581),
            product_re_out=>mul_re_out(581),
            product_im_out=>mul_im_out(581)
        );

    UMUL_582 : complex_multiplier
    generic map(
            re_multiplicator=>15492, --- 0.945556640625 + j-0.325256347656
            im_multiplicator=>-5329
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(582),
            data_im_in=>first_stage_im_out(582),
            product_re_out=>mul_re_out(582),
            product_im_out=>mul_im_out(582)
        );

    UMUL_583 : complex_multiplier
    generic map(
            re_multiplicator=>15175, --- 0.926208496094 + j-0.376953125
            im_multiplicator=>-6176
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(583),
            data_im_in=>first_stage_im_out(583),
            product_re_out=>mul_re_out(583),
            product_im_out=>mul_im_out(583)
        );

    UMUL_584 : complex_multiplier
    generic map(
            re_multiplicator=>14810, --- 0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(584),
            data_im_in=>first_stage_im_out(584),
            product_re_out=>mul_re_out(584),
            product_im_out=>mul_im_out(584)
        );

    UMUL_585 : complex_multiplier
    generic map(
            re_multiplicator=>14401, --- 0.878967285156 + j-0.476745605469
            im_multiplicator=>-7811
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(585),
            data_im_in=>first_stage_im_out(585),
            product_re_out=>mul_re_out(585),
            product_im_out=>mul_im_out(585)
        );

    UMUL_586 : complex_multiplier
    generic map(
            re_multiplicator=>13948, --- 0.851318359375 + j-0.524536132812
            im_multiplicator=>-8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(586),
            data_im_in=>first_stage_im_out(586),
            product_re_out=>mul_re_out(586),
            product_im_out=>mul_im_out(586)
        );

    UMUL_587 : complex_multiplier
    generic map(
            re_multiplicator=>13452, --- 0.821044921875 + j-0.570739746094
            im_multiplicator=>-9351
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(587),
            data_im_in=>first_stage_im_out(587),
            product_re_out=>mul_re_out(587),
            product_im_out=>mul_im_out(587)
        );

    UMUL_588 : complex_multiplier
    generic map(
            re_multiplicator=>12916, --- 0.788330078125 + j-0.615173339844
            im_multiplicator=>-10079
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(588),
            data_im_in=>first_stage_im_out(588),
            product_re_out=>mul_re_out(588),
            product_im_out=>mul_im_out(588)
        );

    UMUL_589 : complex_multiplier
    generic map(
            re_multiplicator=>12340, --- 0.753173828125 + j-0.657775878906
            im_multiplicator=>-10777
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(589),
            data_im_in=>first_stage_im_out(589),
            product_re_out=>mul_re_out(589),
            product_im_out=>mul_im_out(589)
        );

    UMUL_590 : complex_multiplier
    generic map(
            re_multiplicator=>11726, --- 0.715698242188 + j-0.698364257812
            im_multiplicator=>-11442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(590),
            data_im_in=>first_stage_im_out(590),
            product_re_out=>mul_re_out(590),
            product_im_out=>mul_im_out(590)
        );

    UMUL_591 : complex_multiplier
    generic map(
            re_multiplicator=>11077, --- 0.676086425781 + j-0.73681640625
            im_multiplicator=>-12072
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(591),
            data_im_in=>first_stage_im_out(591),
            product_re_out=>mul_re_out(591),
            product_im_out=>mul_im_out(591)
        );

    UMUL_592 : complex_multiplier
    generic map(
            re_multiplicator=>10393, --- 0.634338378906 + j-0.773010253906
            im_multiplicator=>-12665
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(592),
            data_im_in=>first_stage_im_out(592),
            product_re_out=>mul_re_out(592),
            product_im_out=>mul_im_out(592)
        );

    UMUL_593 : complex_multiplier
    generic map(
            re_multiplicator=>9679, --- 0.590759277344 + j-0.806823730469
            im_multiplicator=>-13219
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(593),
            data_im_in=>first_stage_im_out(593),
            product_re_out=>mul_re_out(593),
            product_im_out=>mul_im_out(593)
        );

    UMUL_594 : complex_multiplier
    generic map(
            re_multiplicator=>8934, --- 0.545288085938 + j-0.838195800781
            im_multiplicator=>-13733
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(594),
            data_im_in=>first_stage_im_out(594),
            product_re_out=>mul_re_out(594),
            product_im_out=>mul_im_out(594)
        );

    UMUL_595 : complex_multiplier
    generic map(
            re_multiplicator=>8162, --- 0.498168945312 + j-0.867004394531
            im_multiplicator=>-14205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(595),
            data_im_in=>first_stage_im_out(595),
            product_re_out=>mul_re_out(595),
            product_im_out=>mul_im_out(595)
        );

    UMUL_596 : complex_multiplier
    generic map(
            re_multiplicator=>7366, --- 0.449584960938 + j-0.893188476562
            im_multiplicator=>-14634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(596),
            data_im_in=>first_stage_im_out(596),
            product_re_out=>mul_re_out(596),
            product_im_out=>mul_im_out(596)
        );

    UMUL_597 : complex_multiplier
    generic map(
            re_multiplicator=>6547, --- 0.399597167969 + j-0.916625976562
            im_multiplicator=>-15018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(597),
            data_im_in=>first_stage_im_out(597),
            product_re_out=>mul_re_out(597),
            product_im_out=>mul_im_out(597)
        );

    UMUL_598 : complex_multiplier
    generic map(
            re_multiplicator=>5708, --- 0.348388671875 + j-0.937316894531
            im_multiplicator=>-15357
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(598),
            data_im_in=>first_stage_im_out(598),
            product_re_out=>mul_re_out(598),
            product_im_out=>mul_im_out(598)
        );

    UMUL_599 : complex_multiplier
    generic map(
            re_multiplicator=>4852, --- 0.296142578125 + j-0.955139160156
            im_multiplicator=>-15649
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(599),
            data_im_in=>first_stage_im_out(599),
            product_re_out=>mul_re_out(599),
            product_im_out=>mul_im_out(599)
        );

    UMUL_600 : complex_multiplier
    generic map(
            re_multiplicator=>3980, --- 0.242919921875 + j-0.969970703125
            im_multiplicator=>-15892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(600),
            data_im_in=>first_stage_im_out(600),
            product_re_out=>mul_re_out(600),
            product_im_out=>mul_im_out(600)
        );

    UMUL_601 : complex_multiplier
    generic map(
            re_multiplicator=>3097, --- 0.189025878906 + j-0.98193359375
            im_multiplicator=>-16088
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(601),
            data_im_in=>first_stage_im_out(601),
            product_re_out=>mul_re_out(601),
            product_im_out=>mul_im_out(601)
        );

    UMUL_602 : complex_multiplier
    generic map(
            re_multiplicator=>2204, --- 0.134521484375 + j-0.990844726562
            im_multiplicator=>-16234
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(602),
            data_im_in=>first_stage_im_out(602),
            product_re_out=>mul_re_out(602),
            product_im_out=>mul_im_out(602)
        );

    UMUL_603 : complex_multiplier
    generic map(
            re_multiplicator=>1305, --- 0.0796508789062 + j-0.996765136719
            im_multiplicator=>-16331
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(603),
            data_im_in=>first_stage_im_out(603),
            product_re_out=>mul_re_out(603),
            product_im_out=>mul_im_out(603)
        );

    UMUL_604 : complex_multiplier
    generic map(
            re_multiplicator=>402, --- 0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(604),
            data_im_in=>first_stage_im_out(604),
            product_re_out=>mul_re_out(604),
            product_im_out=>mul_im_out(604)
        );

    UMUL_605 : complex_multiplier
    generic map(
            re_multiplicator=>-502, --- -0.0306396484375 + j-0.99951171875
            im_multiplicator=>-16376
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(605),
            data_im_in=>first_stage_im_out(605),
            product_re_out=>mul_re_out(605),
            product_im_out=>mul_im_out(605)
        );

    UMUL_606 : complex_multiplier
    generic map(
            re_multiplicator=>-1405, --- -0.0857543945312 + j-0.996276855469
            im_multiplicator=>-16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(606),
            data_im_in=>first_stage_im_out(606),
            product_re_out=>mul_re_out(606),
            product_im_out=>mul_im_out(606)
        );

    UMUL_607 : complex_multiplier
    generic map(
            re_multiplicator=>-2304, --- -0.140625 + j-0.990051269531
            im_multiplicator=>-16221
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(607),
            data_im_in=>first_stage_im_out(607),
            product_re_out=>mul_re_out(607),
            product_im_out=>mul_im_out(607)
        );

    UDELAY_608_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(608),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(608)
        );
    UDELAY_608_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(608),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(608)
        );
    USHIFTER_608_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(608),
            data_out=>mul_re_out(608)
        );
    USHIFTER_608_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(608),
            data_out=>mul_im_out(608)
        );

    UMUL_609 : complex_multiplier
    generic map(
            re_multiplicator=>16356, --- 0.998291015625 + j-0.0582275390625
            im_multiplicator=>-954
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(609),
            data_im_in=>first_stage_im_out(609),
            product_re_out=>mul_re_out(609),
            product_im_out=>mul_im_out(609)
        );

    UMUL_610 : complex_multiplier
    generic map(
            re_multiplicator=>16272, --- 0.9931640625 + j-0.116271972656
            im_multiplicator=>-1905
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(610),
            data_im_in=>first_stage_im_out(610),
            product_re_out=>mul_re_out(610),
            product_im_out=>mul_im_out(610)
        );

    UMUL_611 : complex_multiplier
    generic map(
            re_multiplicator=>16134, --- 0.984741210938 + j-0.173950195312
            im_multiplicator=>-2850
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(611),
            data_im_in=>first_stage_im_out(611),
            product_re_out=>mul_re_out(611),
            product_im_out=>mul_im_out(611)
        );

    UMUL_612 : complex_multiplier
    generic map(
            re_multiplicator=>15940, --- 0.972900390625 + j-0.231018066406
            im_multiplicator=>-3785
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(612),
            data_im_in=>first_stage_im_out(612),
            product_re_out=>mul_re_out(612),
            product_im_out=>mul_im_out(612)
        );

    UMUL_613 : complex_multiplier
    generic map(
            re_multiplicator=>15693, --- 0.957824707031 + j-0.287292480469
            im_multiplicator=>-4707
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(613),
            data_im_in=>first_stage_im_out(613),
            product_re_out=>mul_re_out(613),
            product_im_out=>mul_im_out(613)
        );

    UMUL_614 : complex_multiplier
    generic map(
            re_multiplicator=>15392, --- 0.939453125 + j-0.342651367188
            im_multiplicator=>-5614
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(614),
            data_im_in=>first_stage_im_out(614),
            product_re_out=>mul_re_out(614),
            product_im_out=>mul_im_out(614)
        );

    UMUL_615 : complex_multiplier
    generic map(
            re_multiplicator=>15038, --- 0.917846679688 + j-0.396789550781
            im_multiplicator=>-6501
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(615),
            data_im_in=>first_stage_im_out(615),
            product_re_out=>mul_re_out(615),
            product_im_out=>mul_im_out(615)
        );

    UMUL_616 : complex_multiplier
    generic map(
            re_multiplicator=>14634, --- 0.893188476562 + j-0.449584960938
            im_multiplicator=>-7366
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(616),
            data_im_in=>first_stage_im_out(616),
            product_re_out=>mul_re_out(616),
            product_im_out=>mul_im_out(616)
        );

    UMUL_617 : complex_multiplier
    generic map(
            re_multiplicator=>14180, --- 0.865478515625 + j-0.500854492188
            im_multiplicator=>-8206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(617),
            data_im_in=>first_stage_im_out(617),
            product_re_out=>mul_re_out(617),
            product_im_out=>mul_im_out(617)
        );

    UMUL_618 : complex_multiplier
    generic map(
            re_multiplicator=>13678, --- 0.834838867188 + j-0.550415039062
            im_multiplicator=>-9018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(618),
            data_im_in=>first_stage_im_out(618),
            product_re_out=>mul_re_out(618),
            product_im_out=>mul_im_out(618)
        );

    UMUL_619 : complex_multiplier
    generic map(
            re_multiplicator=>13129, --- 0.801330566406 + j-0.59814453125
            im_multiplicator=>-9800
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(619),
            data_im_in=>first_stage_im_out(619),
            product_re_out=>mul_re_out(619),
            product_im_out=>mul_im_out(619)
        );

    UMUL_620 : complex_multiplier
    generic map(
            re_multiplicator=>12536, --- 0.76513671875 + j-0.643798828125
            im_multiplicator=>-10548
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(620),
            data_im_in=>first_stage_im_out(620),
            product_re_out=>mul_re_out(620),
            product_im_out=>mul_im_out(620)
        );

    UMUL_621 : complex_multiplier
    generic map(
            re_multiplicator=>11900, --- 0.726318359375 + j-0.687255859375
            im_multiplicator=>-11260
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(621),
            data_im_in=>first_stage_im_out(621),
            product_re_out=>mul_re_out(621),
            product_im_out=>mul_im_out(621)
        );

    UMUL_622 : complex_multiplier
    generic map(
            re_multiplicator=>11224, --- 0.68505859375 + j-0.728454589844
            im_multiplicator=>-11935
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(622),
            data_im_in=>first_stage_im_out(622),
            product_re_out=>mul_re_out(622),
            product_im_out=>mul_im_out(622)
        );

    UMUL_623 : complex_multiplier
    generic map(
            re_multiplicator=>10510, --- 0.641479492188 + j-0.76708984375
            im_multiplicator=>-12568
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(623),
            data_im_in=>first_stage_im_out(623),
            product_re_out=>mul_re_out(623),
            product_im_out=>mul_im_out(623)
        );

    UMUL_624 : complex_multiplier
    generic map(
            re_multiplicator=>9759, --- 0.595642089844 + j-0.803161621094
            im_multiplicator=>-13159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(624),
            data_im_in=>first_stage_im_out(624),
            product_re_out=>mul_re_out(624),
            product_im_out=>mul_im_out(624)
        );

    UMUL_625 : complex_multiplier
    generic map(
            re_multiplicator=>8976, --- 0.5478515625 + j-0.836486816406
            im_multiplicator=>-13705
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(625),
            data_im_in=>first_stage_im_out(625),
            product_re_out=>mul_re_out(625),
            product_im_out=>mul_im_out(625)
        );

    UMUL_626 : complex_multiplier
    generic map(
            re_multiplicator=>8162, --- 0.498168945312 + j-0.867004394531
            im_multiplicator=>-14205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(626),
            data_im_in=>first_stage_im_out(626),
            product_re_out=>mul_re_out(626),
            product_im_out=>mul_im_out(626)
        );

    UMUL_627 : complex_multiplier
    generic map(
            re_multiplicator=>7321, --- 0.446838378906 + j-0.894592285156
            im_multiplicator=>-14657
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(627),
            data_im_in=>first_stage_im_out(627),
            product_re_out=>mul_re_out(627),
            product_im_out=>mul_im_out(627)
        );

    UMUL_628 : complex_multiplier
    generic map(
            re_multiplicator=>6455, --- 0.393981933594 + j-0.919067382812
            im_multiplicator=>-15058
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(628),
            data_im_in=>first_stage_im_out(628),
            product_re_out=>mul_re_out(628),
            product_im_out=>mul_im_out(628)
        );

    UMUL_629 : complex_multiplier
    generic map(
            re_multiplicator=>5566, --- 0.339721679688 + j-0.940490722656
            im_multiplicator=>-15409
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(629),
            data_im_in=>first_stage_im_out(629),
            product_re_out=>mul_re_out(629),
            product_im_out=>mul_im_out(629)
        );

    UMUL_630 : complex_multiplier
    generic map(
            re_multiplicator=>4659, --- 0.284362792969 + j-0.958679199219
            im_multiplicator=>-15707
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(630),
            data_im_in=>first_stage_im_out(630),
            product_re_out=>mul_re_out(630),
            product_im_out=>mul_im_out(630)
        );

    UMUL_631 : complex_multiplier
    generic map(
            re_multiplicator=>3736, --- 0.22802734375 + j-0.9736328125
            im_multiplicator=>-15952
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(631),
            data_im_in=>first_stage_im_out(631),
            product_re_out=>mul_re_out(631),
            product_im_out=>mul_im_out(631)
        );

    UMUL_632 : complex_multiplier
    generic map(
            re_multiplicator=>2801, --- 0.170959472656 + j-0.985229492188
            im_multiplicator=>-16142
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(632),
            data_im_in=>first_stage_im_out(632),
            product_re_out=>mul_re_out(632),
            product_im_out=>mul_im_out(632)
        );

    UMUL_633 : complex_multiplier
    generic map(
            re_multiplicator=>1855, --- 0.113220214844 + j-0.993530273438
            im_multiplicator=>-16278
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(633),
            data_im_in=>first_stage_im_out(633),
            product_re_out=>mul_re_out(633),
            product_im_out=>mul_im_out(633)
        );

    UMUL_634 : complex_multiplier
    generic map(
            re_multiplicator=>904, --- 0.05517578125 + j-0.998474121094
            im_multiplicator=>-16359
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(634),
            data_im_in=>first_stage_im_out(634),
            product_re_out=>mul_re_out(634),
            product_im_out=>mul_im_out(634)
        );

    UMUL_635 : complex_multiplier
    generic map(
            re_multiplicator=>-50, --- -0.0030517578125 + j-0.999938964844
            im_multiplicator=>-16383
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(635),
            data_im_in=>first_stage_im_out(635),
            product_re_out=>mul_re_out(635),
            product_im_out=>mul_im_out(635)
        );

    UMUL_636 : complex_multiplier
    generic map(
            re_multiplicator=>-1004, --- -0.061279296875 + j-0.998107910156
            im_multiplicator=>-16353
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(636),
            data_im_in=>first_stage_im_out(636),
            product_re_out=>mul_re_out(636),
            product_im_out=>mul_im_out(636)
        );

    UMUL_637 : complex_multiplier
    generic map(
            re_multiplicator=>-1955, --- -0.119323730469 + j-0.992797851562
            im_multiplicator=>-16266
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(637),
            data_im_in=>first_stage_im_out(637),
            product_re_out=>mul_re_out(637),
            product_im_out=>mul_im_out(637)
        );

    UMUL_638 : complex_multiplier
    generic map(
            re_multiplicator=>-2900, --- -0.177001953125 + j-0.984191894531
            im_multiplicator=>-16125
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(638),
            data_im_in=>first_stage_im_out(638),
            product_re_out=>mul_re_out(638),
            product_im_out=>mul_im_out(638)
        );

    UMUL_639 : complex_multiplier
    generic map(
            re_multiplicator=>-3834, --- -0.234008789062 + j-0.97216796875
            im_multiplicator=>-15928
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(639),
            data_im_in=>first_stage_im_out(639),
            product_re_out=>mul_re_out(639),
            product_im_out=>mul_im_out(639)
        );

    UDELAY_640_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(640),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(640)
        );
    UDELAY_640_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(640),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(640)
        );
    USHIFTER_640_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(640),
            data_out=>mul_re_out(640)
        );
    USHIFTER_640_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(640),
            data_out=>mul_im_out(640)
        );

    UMUL_641 : complex_multiplier
    generic map(
            re_multiplicator=>16353, --- 0.998107910156 + j-0.061279296875
            im_multiplicator=>-1004
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(641),
            data_im_in=>first_stage_im_out(641),
            product_re_out=>mul_re_out(641),
            product_im_out=>mul_im_out(641)
        );

    UMUL_642 : complex_multiplier
    generic map(
            re_multiplicator=>16260, --- 0.992431640625 + j-0.122375488281
            im_multiplicator=>-2005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(642),
            data_im_in=>first_stage_im_out(642),
            product_re_out=>mul_re_out(642),
            product_im_out=>mul_im_out(642)
        );

    UMUL_643 : complex_multiplier
    generic map(
            re_multiplicator=>16107, --- 0.983093261719 + j-0.182983398438
            im_multiplicator=>-2998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(643),
            data_im_in=>first_stage_im_out(643),
            product_re_out=>mul_re_out(643),
            product_im_out=>mul_im_out(643)
        );

    UMUL_644 : complex_multiplier
    generic map(
            re_multiplicator=>15892, --- 0.969970703125 + j-0.242919921875
            im_multiplicator=>-3980
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(644),
            data_im_in=>first_stage_im_out(644),
            product_re_out=>mul_re_out(644),
            product_im_out=>mul_im_out(644)
        );

    UMUL_645 : complex_multiplier
    generic map(
            re_multiplicator=>15618, --- 0.953247070312 + j-0.302001953125
            im_multiplicator=>-4948
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(645),
            data_im_in=>first_stage_im_out(645),
            product_re_out=>mul_re_out(645),
            product_im_out=>mul_im_out(645)
        );

    UMUL_646 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(646),
            data_im_in=>first_stage_im_out(646),
            product_re_out=>mul_re_out(646),
            product_im_out=>mul_im_out(646)
        );

    UMUL_647 : complex_multiplier
    generic map(
            re_multiplicator=>14895, --- 0.909118652344 + j-0.416381835938
            im_multiplicator=>-6822
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(647),
            data_im_in=>first_stage_im_out(647),
            product_re_out=>mul_re_out(647),
            product_im_out=>mul_im_out(647)
        );

    UMUL_648 : complex_multiplier
    generic map(
            re_multiplicator=>14449, --- 0.881896972656 + j-0.471374511719
            im_multiplicator=>-7723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(648),
            data_im_in=>first_stage_im_out(648),
            product_re_out=>mul_re_out(648),
            product_im_out=>mul_im_out(648)
        );

    UMUL_649 : complex_multiplier
    generic map(
            re_multiplicator=>13948, --- 0.851318359375 + j-0.524536132812
            im_multiplicator=>-8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(649),
            data_im_in=>first_stage_im_out(649),
            product_re_out=>mul_re_out(649),
            product_im_out=>mul_im_out(649)
        );

    UMUL_650 : complex_multiplier
    generic map(
            re_multiplicator=>13395, --- 0.817565917969 + j-0.575805664062
            im_multiplicator=>-9434
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(650),
            data_im_in=>first_stage_im_out(650),
            product_re_out=>mul_re_out(650),
            product_im_out=>mul_im_out(650)
        );

    UMUL_651 : complex_multiplier
    generic map(
            re_multiplicator=>12791, --- 0.780700683594 + j-0.624816894531
            im_multiplicator=>-10237
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(651),
            data_im_in=>first_stage_im_out(651),
            product_re_out=>mul_re_out(651),
            product_im_out=>mul_im_out(651)
        );

    UMUL_652 : complex_multiplier
    generic map(
            re_multiplicator=>12139, --- 0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(652),
            data_im_in=>first_stage_im_out(652),
            product_re_out=>mul_re_out(652),
            product_im_out=>mul_im_out(652)
        );

    UMUL_653 : complex_multiplier
    generic map(
            re_multiplicator=>11442, --- 0.698364257812 + j-0.715698242188
            im_multiplicator=>-11726
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(653),
            data_im_in=>first_stage_im_out(653),
            product_re_out=>mul_re_out(653),
            product_im_out=>mul_im_out(653)
        );

    UMUL_654 : complex_multiplier
    generic map(
            re_multiplicator=>10701, --- 0.653137207031 + j-0.757202148438
            im_multiplicator=>-12406
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(654),
            data_im_in=>first_stage_im_out(654),
            product_re_out=>mul_re_out(654),
            product_im_out=>mul_im_out(654)
        );

    UMUL_655 : complex_multiplier
    generic map(
            re_multiplicator=>9920, --- 0.60546875 + j-0.795776367188
            im_multiplicator=>-13038
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(655),
            data_im_in=>first_stage_im_out(655),
            product_re_out=>mul_re_out(655),
            product_im_out=>mul_im_out(655)
        );

    UMUL_656 : complex_multiplier
    generic map(
            re_multiplicator=>9102, --- 0.555541992188 + j-0.831420898438
            im_multiplicator=>-13622
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(656),
            data_im_in=>first_stage_im_out(656),
            product_re_out=>mul_re_out(656),
            product_im_out=>mul_im_out(656)
        );

    UMUL_657 : complex_multiplier
    generic map(
            re_multiplicator=>8249, --- 0.503479003906 + j-0.863952636719
            im_multiplicator=>-14155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(657),
            data_im_in=>first_stage_im_out(657),
            product_re_out=>mul_re_out(657),
            product_im_out=>mul_im_out(657)
        );

    UMUL_658 : complex_multiplier
    generic map(
            re_multiplicator=>7366, --- 0.449584960938 + j-0.893188476562
            im_multiplicator=>-14634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(658),
            data_im_in=>first_stage_im_out(658),
            product_re_out=>mul_re_out(658),
            product_im_out=>mul_im_out(658)
        );

    UMUL_659 : complex_multiplier
    generic map(
            re_multiplicator=>6455, --- 0.393981933594 + j-0.919067382812
            im_multiplicator=>-15058
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(659),
            data_im_in=>first_stage_im_out(659),
            product_re_out=>mul_re_out(659),
            product_im_out=>mul_im_out(659)
        );

    UMUL_660 : complex_multiplier
    generic map(
            re_multiplicator=>5519, --- 0.336853027344 + j-0.941528320312
            im_multiplicator=>-15426
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(660),
            data_im_in=>first_stage_im_out(660),
            product_re_out=>mul_re_out(660),
            product_im_out=>mul_im_out(660)
        );

    UMUL_661 : complex_multiplier
    generic map(
            re_multiplicator=>4563, --- 0.278503417969 + j-0.960388183594
            im_multiplicator=>-15735
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(661),
            data_im_in=>first_stage_im_out(661),
            product_re_out=>mul_re_out(661),
            product_im_out=>mul_im_out(661)
        );

    UMUL_662 : complex_multiplier
    generic map(
            re_multiplicator=>3589, --- 0.219055175781 + j-0.975646972656
            im_multiplicator=>-15985
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(662),
            data_im_in=>first_stage_im_out(662),
            product_re_out=>mul_re_out(662),
            product_im_out=>mul_im_out(662)
        );

    UMUL_663 : complex_multiplier
    generic map(
            re_multiplicator=>2602, --- 0.158813476562 + j-0.987243652344
            im_multiplicator=>-16175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(663),
            data_im_in=>first_stage_im_out(663),
            product_re_out=>mul_re_out(663),
            product_im_out=>mul_im_out(663)
        );

    UMUL_664 : complex_multiplier
    generic map(
            re_multiplicator=>1605, --- 0.0979614257812 + j-0.995178222656
            im_multiplicator=>-16305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(664),
            data_im_in=>first_stage_im_out(664),
            product_re_out=>mul_re_out(664),
            product_im_out=>mul_im_out(664)
        );

    UMUL_665 : complex_multiplier
    generic map(
            re_multiplicator=>603, --- 0.0368041992188 + j-0.999267578125
            im_multiplicator=>-16372
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(665),
            data_im_in=>first_stage_im_out(665),
            product_re_out=>mul_re_out(665),
            product_im_out=>mul_im_out(665)
        );

    UMUL_666 : complex_multiplier
    generic map(
            re_multiplicator=>-402, --- -0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(666),
            data_im_in=>first_stage_im_out(666),
            product_re_out=>mul_re_out(666),
            product_im_out=>mul_im_out(666)
        );

    UMUL_667 : complex_multiplier
    generic map(
            re_multiplicator=>-1405, --- -0.0857543945312 + j-0.996276855469
            im_multiplicator=>-16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(667),
            data_im_in=>first_stage_im_out(667),
            product_re_out=>mul_re_out(667),
            product_im_out=>mul_im_out(667)
        );

    UMUL_668 : complex_multiplier
    generic map(
            re_multiplicator=>-2404, --- -0.146728515625 + j-0.989135742188
            im_multiplicator=>-16206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(668),
            data_im_in=>first_stage_im_out(668),
            product_re_out=>mul_re_out(668),
            product_im_out=>mul_im_out(668)
        );

    UMUL_669 : complex_multiplier
    generic map(
            re_multiplicator=>-3393, --- -0.207092285156 + j-0.978271484375
            im_multiplicator=>-16028
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(669),
            data_im_in=>first_stage_im_out(669),
            product_re_out=>mul_re_out(669),
            product_im_out=>mul_im_out(669)
        );

    UMUL_670 : complex_multiplier
    generic map(
            re_multiplicator=>-4369, --- -0.266662597656 + j-0.963745117188
            im_multiplicator=>-15790
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(670),
            data_im_in=>first_stage_im_out(670),
            product_re_out=>mul_re_out(670),
            product_im_out=>mul_im_out(670)
        );

    UMUL_671 : complex_multiplier
    generic map(
            re_multiplicator=>-5329, --- -0.325256347656 + j-0.945556640625
            im_multiplicator=>-15492
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(671),
            data_im_in=>first_stage_im_out(671),
            product_re_out=>mul_re_out(671),
            product_im_out=>mul_im_out(671)
        );

    UDELAY_672_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(672),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(672)
        );
    UDELAY_672_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(672),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(672)
        );
    USHIFTER_672_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(672),
            data_out=>mul_re_out(672)
        );
    USHIFTER_672_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(672),
            data_out=>mul_im_out(672)
        );

    UMUL_673 : complex_multiplier
    generic map(
            re_multiplicator=>16350, --- 0.997924804688 + j-0.0643310546875
            im_multiplicator=>-1054
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(673),
            data_im_in=>first_stage_im_out(673),
            product_re_out=>mul_re_out(673),
            product_im_out=>mul_im_out(673)
        );

    UMUL_674 : complex_multiplier
    generic map(
            re_multiplicator=>16248, --- 0.99169921875 + j-0.128479003906
            im_multiplicator=>-2105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(674),
            data_im_in=>first_stage_im_out(674),
            product_re_out=>mul_re_out(674),
            product_im_out=>mul_im_out(674)
        );

    UMUL_675 : complex_multiplier
    generic map(
            re_multiplicator=>16078, --- 0.981323242188 + j-0.192077636719
            im_multiplicator=>-3147
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(675),
            data_im_in=>first_stage_im_out(675),
            product_re_out=>mul_re_out(675),
            product_im_out=>mul_im_out(675)
        );

    UMUL_676 : complex_multiplier
    generic map(
            re_multiplicator=>15842, --- 0.966918945312 + j-0.254821777344
            im_multiplicator=>-4175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(676),
            data_im_in=>first_stage_im_out(676),
            product_re_out=>mul_re_out(676),
            product_im_out=>mul_im_out(676)
        );

    UMUL_677 : complex_multiplier
    generic map(
            re_multiplicator=>15541, --- 0.948547363281 + j-0.316589355469
            im_multiplicator=>-5187
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(677),
            data_im_in=>first_stage_im_out(677),
            product_re_out=>mul_re_out(677),
            product_im_out=>mul_im_out(677)
        );

    UMUL_678 : complex_multiplier
    generic map(
            re_multiplicator=>15175, --- 0.926208496094 + j-0.376953125
            im_multiplicator=>-6176
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(678),
            data_im_in=>first_stage_im_out(678),
            product_re_out=>mul_re_out(678),
            product_im_out=>mul_im_out(678)
        );

    UMUL_679 : complex_multiplier
    generic map(
            re_multiplicator=>14745, --- 0.899963378906 + j-0.435852050781
            im_multiplicator=>-7141
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(679),
            data_im_in=>first_stage_im_out(679),
            product_re_out=>mul_re_out(679),
            product_im_out=>mul_im_out(679)
        );

    UMUL_680 : complex_multiplier
    generic map(
            re_multiplicator=>14255, --- 0.870056152344 + j-0.492858886719
            im_multiplicator=>-8075
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(680),
            data_im_in=>first_stage_im_out(680),
            product_re_out=>mul_re_out(680),
            product_im_out=>mul_im_out(680)
        );

    UMUL_681 : complex_multiplier
    generic map(
            re_multiplicator=>13705, --- 0.836486816406 + j-0.5478515625
            im_multiplicator=>-8976
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(681),
            data_im_in=>first_stage_im_out(681),
            product_re_out=>mul_re_out(681),
            product_im_out=>mul_im_out(681)
        );

    UMUL_682 : complex_multiplier
    generic map(
            re_multiplicator=>13099, --- 0.799499511719 + j-0.6005859375
            im_multiplicator=>-9840
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(682),
            data_im_in=>first_stage_im_out(682),
            product_re_out=>mul_re_out(682),
            product_im_out=>mul_im_out(682)
        );

    UMUL_683 : complex_multiplier
    generic map(
            re_multiplicator=>12438, --- 0.759155273438 + j-0.650817871094
            im_multiplicator=>-10663
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(683),
            data_im_in=>first_stage_im_out(683),
            product_re_out=>mul_re_out(683),
            product_im_out=>mul_im_out(683)
        );

    UMUL_684 : complex_multiplier
    generic map(
            re_multiplicator=>11726, --- 0.715698242188 + j-0.698364257812
            im_multiplicator=>-11442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(684),
            data_im_in=>first_stage_im_out(684),
            product_re_out=>mul_re_out(684),
            product_im_out=>mul_im_out(684)
        );

    UMUL_685 : complex_multiplier
    generic map(
            re_multiplicator=>10965, --- 0.669250488281 + j-0.742980957031
            im_multiplicator=>-12173
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(685),
            data_im_in=>first_stage_im_out(685),
            product_re_out=>mul_re_out(685),
            product_im_out=>mul_im_out(685)
        );

    UMUL_686 : complex_multiplier
    generic map(
            re_multiplicator=>10159, --- 0.620056152344 + j-0.784545898438
            im_multiplicator=>-12854
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(686),
            data_im_in=>first_stage_im_out(686),
            product_re_out=>mul_re_out(686),
            product_im_out=>mul_im_out(686)
        );

    UMUL_687 : complex_multiplier
    generic map(
            re_multiplicator=>9310, --- 0.568237304688 + j-0.822814941406
            im_multiplicator=>-13481
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(687),
            data_im_in=>first_stage_im_out(687),
            product_re_out=>mul_re_out(687),
            product_im_out=>mul_im_out(687)
        );

    UMUL_688 : complex_multiplier
    generic map(
            re_multiplicator=>8423, --- 0.514099121094 + j-0.857727050781
            im_multiplicator=>-14053
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(688),
            data_im_in=>first_stage_im_out(688),
            product_re_out=>mul_re_out(688),
            product_im_out=>mul_im_out(688)
        );

    UMUL_689 : complex_multiplier
    generic map(
            re_multiplicator=>7500, --- 0.457763671875 + j-0.889038085938
            im_multiplicator=>-14566
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(689),
            data_im_in=>first_stage_im_out(689),
            product_re_out=>mul_re_out(689),
            product_im_out=>mul_im_out(689)
        );

    UMUL_690 : complex_multiplier
    generic map(
            re_multiplicator=>6547, --- 0.399597167969 + j-0.916625976562
            im_multiplicator=>-15018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(690),
            data_im_in=>first_stage_im_out(690),
            product_re_out=>mul_re_out(690),
            product_im_out=>mul_im_out(690)
        );

    UMUL_691 : complex_multiplier
    generic map(
            re_multiplicator=>5566, --- 0.339721679688 + j-0.940490722656
            im_multiplicator=>-15409
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(691),
            data_im_in=>first_stage_im_out(691),
            product_re_out=>mul_re_out(691),
            product_im_out=>mul_im_out(691)
        );

    UMUL_692 : complex_multiplier
    generic map(
            re_multiplicator=>4563, --- 0.278503417969 + j-0.960388183594
            im_multiplicator=>-15735
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(692),
            data_im_in=>first_stage_im_out(692),
            product_re_out=>mul_re_out(692),
            product_im_out=>mul_im_out(692)
        );

    UMUL_693 : complex_multiplier
    generic map(
            re_multiplicator=>3540, --- 0.216064453125 + j-0.976318359375
            im_multiplicator=>-15996
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(693),
            data_im_in=>first_stage_im_out(693),
            product_re_out=>mul_re_out(693),
            product_im_out=>mul_im_out(693)
        );

    UMUL_694 : complex_multiplier
    generic map(
            re_multiplicator=>2503, --- 0.152770996094 + j-0.988220214844
            im_multiplicator=>-16191
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(694),
            data_im_in=>first_stage_im_out(694),
            product_re_out=>mul_re_out(694),
            product_im_out=>mul_im_out(694)
        );

    UMUL_695 : complex_multiplier
    generic map(
            re_multiplicator=>1455, --- 0.0888061523438 + j-0.996032714844
            im_multiplicator=>-16319
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(695),
            data_im_in=>first_stage_im_out(695),
            product_re_out=>mul_re_out(695),
            product_im_out=>mul_im_out(695)
        );

    UMUL_696 : complex_multiplier
    generic map(
            re_multiplicator=>402, --- 0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(696),
            data_im_in=>first_stage_im_out(696),
            product_re_out=>mul_re_out(696),
            product_im_out=>mul_im_out(696)
        );

    UMUL_697 : complex_multiplier
    generic map(
            re_multiplicator=>-653, --- -0.0398559570312 + j-0.999145507812
            im_multiplicator=>-16370
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(697),
            data_im_in=>first_stage_im_out(697),
            product_re_out=>mul_re_out(697),
            product_im_out=>mul_im_out(697)
        );

    UMUL_698 : complex_multiplier
    generic map(
            re_multiplicator=>-1705, --- -0.104064941406 + j-0.994506835938
            im_multiplicator=>-16294
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(698),
            data_im_in=>first_stage_im_out(698),
            product_re_out=>mul_re_out(698),
            product_im_out=>mul_im_out(698)
        );

    UMUL_699 : complex_multiplier
    generic map(
            re_multiplicator=>-2751, --- -0.167907714844 + j-0.985778808594
            im_multiplicator=>-16151
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(699),
            data_im_in=>first_stage_im_out(699),
            product_re_out=>mul_re_out(699),
            product_im_out=>mul_im_out(699)
        );

    UMUL_700 : complex_multiplier
    generic map(
            re_multiplicator=>-3785, --- -0.231018066406 + j-0.972900390625
            im_multiplicator=>-15940
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(700),
            data_im_in=>first_stage_im_out(700),
            product_re_out=>mul_re_out(700),
            product_im_out=>mul_im_out(700)
        );

    UMUL_701 : complex_multiplier
    generic map(
            re_multiplicator=>-4804, --- -0.293212890625 + j-0.955993652344
            im_multiplicator=>-15663
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(701),
            data_im_in=>first_stage_im_out(701),
            product_re_out=>mul_re_out(701),
            product_im_out=>mul_im_out(701)
        );

    UMUL_702 : complex_multiplier
    generic map(
            re_multiplicator=>-5802, --- -0.354125976562 + j-0.935180664062
            im_multiplicator=>-15322
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(702),
            data_im_in=>first_stage_im_out(702),
            product_re_out=>mul_re_out(702),
            product_im_out=>mul_im_out(702)
        );

    UMUL_703 : complex_multiplier
    generic map(
            re_multiplicator=>-6777, --- -0.413635253906 + j-0.910400390625
            im_multiplicator=>-14916
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(703),
            data_im_in=>first_stage_im_out(703),
            product_re_out=>mul_re_out(703),
            product_im_out=>mul_im_out(703)
        );

    UDELAY_704_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(704),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(704)
        );
    UDELAY_704_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(704),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(704)
        );
    USHIFTER_704_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(704),
            data_out=>mul_re_out(704)
        );
    USHIFTER_704_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(704),
            data_out=>mul_im_out(704)
        );

    UMUL_705 : complex_multiplier
    generic map(
            re_multiplicator=>16346, --- 0.997680664062 + j-0.0674438476562
            im_multiplicator=>-1105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(705),
            data_im_in=>first_stage_im_out(705),
            product_re_out=>mul_re_out(705),
            product_im_out=>mul_im_out(705)
        );

    UMUL_706 : complex_multiplier
    generic map(
            re_multiplicator=>16234, --- 0.990844726562 + j-0.134521484375
            im_multiplicator=>-2204
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(706),
            data_im_in=>first_stage_im_out(706),
            product_re_out=>mul_re_out(706),
            product_im_out=>mul_im_out(706)
        );

    UMUL_707 : complex_multiplier
    generic map(
            re_multiplicator=>16049, --- 0.979553222656 + j-0.201049804688
            im_multiplicator=>-3294
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(707),
            data_im_in=>first_stage_im_out(707),
            product_re_out=>mul_re_out(707),
            product_im_out=>mul_im_out(707)
        );

    UMUL_708 : complex_multiplier
    generic map(
            re_multiplicator=>15790, --- 0.963745117188 + j-0.266662597656
            im_multiplicator=>-4369
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(708),
            data_im_in=>first_stage_im_out(708),
            product_re_out=>mul_re_out(708),
            product_im_out=>mul_im_out(708)
        );

    UMUL_709 : complex_multiplier
    generic map(
            re_multiplicator=>15459, --- 0.943542480469 + j-0.3310546875
            im_multiplicator=>-5424
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(709),
            data_im_in=>first_stage_im_out(709),
            product_re_out=>mul_re_out(709),
            product_im_out=>mul_im_out(709)
        );

    UMUL_710 : complex_multiplier
    generic map(
            re_multiplicator=>15058, --- 0.919067382812 + j-0.393981933594
            im_multiplicator=>-6455
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(710),
            data_im_in=>first_stage_im_out(710),
            product_re_out=>mul_re_out(710),
            product_im_out=>mul_im_out(710)
        );

    UMUL_711 : complex_multiplier
    generic map(
            re_multiplicator=>14589, --- 0.890441894531 + j-0.455078125
            im_multiplicator=>-7456
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(711),
            data_im_in=>first_stage_im_out(711),
            product_re_out=>mul_re_out(711),
            product_im_out=>mul_im_out(711)
        );

    UMUL_712 : complex_multiplier
    generic map(
            re_multiplicator=>14053, --- 0.857727050781 + j-0.514099121094
            im_multiplicator=>-8423
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(712),
            data_im_in=>first_stage_im_out(712),
            product_re_out=>mul_re_out(712),
            product_im_out=>mul_im_out(712)
        );

    UMUL_713 : complex_multiplier
    generic map(
            re_multiplicator=>13452, --- 0.821044921875 + j-0.570739746094
            im_multiplicator=>-9351
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(713),
            data_im_in=>first_stage_im_out(713),
            product_re_out=>mul_re_out(713),
            product_im_out=>mul_im_out(713)
        );

    UMUL_714 : complex_multiplier
    generic map(
            re_multiplicator=>12791, --- 0.780700683594 + j-0.624816894531
            im_multiplicator=>-10237
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(714),
            data_im_in=>first_stage_im_out(714),
            product_re_out=>mul_re_out(714),
            product_im_out=>mul_im_out(714)
        );

    UMUL_715 : complex_multiplier
    generic map(
            re_multiplicator=>12072, --- 0.73681640625 + j-0.676086425781
            im_multiplicator=>-11077
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(715),
            data_im_in=>first_stage_im_out(715),
            product_re_out=>mul_re_out(715),
            product_im_out=>mul_im_out(715)
        );

    UMUL_716 : complex_multiplier
    generic map(
            re_multiplicator=>11297, --- 0.689514160156 + j-0.724243164062
            im_multiplicator=>-11866
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(716),
            data_im_in=>first_stage_im_out(716),
            product_re_out=>mul_re_out(716),
            product_im_out=>mul_im_out(716)
        );

    UMUL_717 : complex_multiplier
    generic map(
            re_multiplicator=>10471, --- 0.639099121094 + j-0.76904296875
            im_multiplicator=>-12600
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(717),
            data_im_in=>first_stage_im_out(717),
            product_re_out=>mul_re_out(717),
            product_im_out=>mul_im_out(717)
        );

    UMUL_718 : complex_multiplier
    generic map(
            re_multiplicator=>9597, --- 0.585754394531 + j-0.810424804688
            im_multiplicator=>-13278
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(718),
            data_im_in=>first_stage_im_out(718),
            product_re_out=>mul_re_out(718),
            product_im_out=>mul_im_out(718)
        );

    UMUL_719 : complex_multiplier
    generic map(
            re_multiplicator=>8680, --- 0.52978515625 + j-0.848083496094
            im_multiplicator=>-13895
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(719),
            data_im_in=>first_stage_im_out(719),
            product_re_out=>mul_re_out(719),
            product_im_out=>mul_im_out(719)
        );

    UMUL_720 : complex_multiplier
    generic map(
            re_multiplicator=>7723, --- 0.471374511719 + j-0.881896972656
            im_multiplicator=>-14449
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(720),
            data_im_in=>first_stage_im_out(720),
            product_re_out=>mul_re_out(720),
            product_im_out=>mul_im_out(720)
        );

    UMUL_721 : complex_multiplier
    generic map(
            re_multiplicator=>6731, --- 0.410827636719 + j-0.911682128906
            im_multiplicator=>-14937
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(721),
            data_im_in=>first_stage_im_out(721),
            product_re_out=>mul_re_out(721),
            product_im_out=>mul_im_out(721)
        );

    UMUL_722 : complex_multiplier
    generic map(
            re_multiplicator=>5708, --- 0.348388671875 + j-0.937316894531
            im_multiplicator=>-15357
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(722),
            data_im_in=>first_stage_im_out(722),
            product_re_out=>mul_re_out(722),
            product_im_out=>mul_im_out(722)
        );

    UMUL_723 : complex_multiplier
    generic map(
            re_multiplicator=>4659, --- 0.284362792969 + j-0.958679199219
            im_multiplicator=>-15707
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(723),
            data_im_in=>first_stage_im_out(723),
            product_re_out=>mul_re_out(723),
            product_im_out=>mul_im_out(723)
        );

    UMUL_724 : complex_multiplier
    generic map(
            re_multiplicator=>3589, --- 0.219055175781 + j-0.975646972656
            im_multiplicator=>-15985
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(724),
            data_im_in=>first_stage_im_out(724),
            product_re_out=>mul_re_out(724),
            product_im_out=>mul_im_out(724)
        );

    UMUL_725 : complex_multiplier
    generic map(
            re_multiplicator=>2503, --- 0.152770996094 + j-0.988220214844
            im_multiplicator=>-16191
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(725),
            data_im_in=>first_stage_im_out(725),
            product_re_out=>mul_re_out(725),
            product_im_out=>mul_im_out(725)
        );

    UMUL_726 : complex_multiplier
    generic map(
            re_multiplicator=>1405, --- 0.0857543945312 + j-0.996276855469
            im_multiplicator=>-16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(726),
            data_im_in=>first_stage_im_out(726),
            product_re_out=>mul_re_out(726),
            product_im_out=>mul_im_out(726)
        );

    UMUL_727 : complex_multiplier
    generic map(
            re_multiplicator=>301, --- 0.0183715820312 + j-0.999816894531
            im_multiplicator=>-16381
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(727),
            data_im_in=>first_stage_im_out(727),
            product_re_out=>mul_re_out(727),
            product_im_out=>mul_im_out(727)
        );

    UMUL_728 : complex_multiplier
    generic map(
            re_multiplicator=>-803, --- -0.0490112304688 + j-0.998779296875
            im_multiplicator=>-16364
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(728),
            data_im_in=>first_stage_im_out(728),
            product_re_out=>mul_re_out(728),
            product_im_out=>mul_im_out(728)
        );

    UMUL_729 : complex_multiplier
    generic map(
            re_multiplicator=>-1905, --- -0.116271972656 + j-0.9931640625
            im_multiplicator=>-16272
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(729),
            data_im_in=>first_stage_im_out(729),
            product_re_out=>mul_re_out(729),
            product_im_out=>mul_im_out(729)
        );

    UMUL_730 : complex_multiplier
    generic map(
            re_multiplicator=>-2998, --- -0.182983398438 + j-0.983093261719
            im_multiplicator=>-16107
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(730),
            data_im_in=>first_stage_im_out(730),
            product_re_out=>mul_re_out(730),
            product_im_out=>mul_im_out(730)
        );

    UMUL_731 : complex_multiplier
    generic map(
            re_multiplicator=>-4078, --- -0.248901367188 + j-0.968505859375
            im_multiplicator=>-15868
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(731),
            data_im_in=>first_stage_im_out(731),
            product_re_out=>mul_re_out(731),
            product_im_out=>mul_im_out(731)
        );

    UMUL_732 : complex_multiplier
    generic map(
            re_multiplicator=>-5139, --- -0.313659667969 + j-0.949523925781
            im_multiplicator=>-15557
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(732),
            data_im_in=>first_stage_im_out(732),
            product_re_out=>mul_re_out(732),
            product_im_out=>mul_im_out(732)
        );

    UMUL_733 : complex_multiplier
    generic map(
            re_multiplicator=>-6176, --- -0.376953125 + j-0.926208496094
            im_multiplicator=>-15175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(733),
            data_im_in=>first_stage_im_out(733),
            product_re_out=>mul_re_out(733),
            product_im_out=>mul_im_out(733)
        );

    UMUL_734 : complex_multiplier
    generic map(
            re_multiplicator=>-7186, --- -0.438598632812 + j-0.898620605469
            im_multiplicator=>-14723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(734),
            data_im_in=>first_stage_im_out(734),
            product_re_out=>mul_re_out(734),
            product_im_out=>mul_im_out(734)
        );

    UMUL_735 : complex_multiplier
    generic map(
            re_multiplicator=>-8162, --- -0.498168945312 + j-0.867004394531
            im_multiplicator=>-14205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(735),
            data_im_in=>first_stage_im_out(735),
            product_re_out=>mul_re_out(735),
            product_im_out=>mul_im_out(735)
        );

    UDELAY_736_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(736),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(736)
        );
    UDELAY_736_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(736),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(736)
        );
    USHIFTER_736_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(736),
            data_out=>mul_re_out(736)
        );
    USHIFTER_736_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(736),
            data_out=>mul_im_out(736)
        );

    UMUL_737 : complex_multiplier
    generic map(
            re_multiplicator=>16343, --- 0.997497558594 + j-0.0704956054688
            im_multiplicator=>-1155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(737),
            data_im_in=>first_stage_im_out(737),
            product_re_out=>mul_re_out(737),
            product_im_out=>mul_im_out(737)
        );

    UMUL_738 : complex_multiplier
    generic map(
            re_multiplicator=>16221, --- 0.990051269531 + j-0.140625
            im_multiplicator=>-2304
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(738),
            data_im_in=>first_stage_im_out(738),
            product_re_out=>mul_re_out(738),
            product_im_out=>mul_im_out(738)
        );

    UMUL_739 : complex_multiplier
    generic map(
            re_multiplicator=>16018, --- 0.977661132812 + j-0.210083007812
            im_multiplicator=>-3442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(739),
            data_im_in=>first_stage_im_out(739),
            product_re_out=>mul_re_out(739),
            product_im_out=>mul_im_out(739)
        );

    UMUL_740 : complex_multiplier
    generic map(
            re_multiplicator=>15735, --- 0.960388183594 + j-0.278503417969
            im_multiplicator=>-4563
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(740),
            data_im_in=>first_stage_im_out(740),
            product_re_out=>mul_re_out(740),
            product_im_out=>mul_im_out(740)
        );

    UMUL_741 : complex_multiplier
    generic map(
            re_multiplicator=>15374, --- 0.938354492188 + j-0.345520019531
            im_multiplicator=>-5661
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(741),
            data_im_in=>first_stage_im_out(741),
            product_re_out=>mul_re_out(741),
            product_im_out=>mul_im_out(741)
        );

    UMUL_742 : complex_multiplier
    generic map(
            re_multiplicator=>14937, --- 0.911682128906 + j-0.410827636719
            im_multiplicator=>-6731
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(742),
            data_im_in=>first_stage_im_out(742),
            product_re_out=>mul_re_out(742),
            product_im_out=>mul_im_out(742)
        );

    UMUL_743 : complex_multiplier
    generic map(
            re_multiplicator=>14425, --- 0.880432128906 + j-0.474060058594
            im_multiplicator=>-7767
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(743),
            data_im_in=>first_stage_im_out(743),
            product_re_out=>mul_re_out(743),
            product_im_out=>mul_im_out(743)
        );

    UMUL_744 : complex_multiplier
    generic map(
            re_multiplicator=>13842, --- 0.844848632812 + j-0.534973144531
            im_multiplicator=>-8765
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(744),
            data_im_in=>first_stage_im_out(744),
            product_re_out=>mul_re_out(744),
            product_im_out=>mul_im_out(744)
        );

    UMUL_745 : complex_multiplier
    generic map(
            re_multiplicator=>13189, --- 0.804992675781 + j-0.593200683594
            im_multiplicator=>-9719
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(745),
            data_im_in=>first_stage_im_out(745),
            product_re_out=>mul_re_out(745),
            product_im_out=>mul_im_out(745)
        );

    UMUL_746 : complex_multiplier
    generic map(
            re_multiplicator=>12471, --- 0.761169433594 + j-0.648498535156
            im_multiplicator=>-10625
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(746),
            data_im_in=>first_stage_im_out(746),
            product_re_out=>mul_re_out(746),
            product_im_out=>mul_im_out(746)
        );

    UMUL_747 : complex_multiplier
    generic map(
            re_multiplicator=>11691, --- 0.713562011719 + j-0.700561523438
            im_multiplicator=>-11478
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(747),
            data_im_in=>first_stage_im_out(747),
            product_re_out=>mul_re_out(747),
            product_im_out=>mul_im_out(747)
        );

    UMUL_748 : complex_multiplier
    generic map(
            re_multiplicator=>10853, --- 0.662414550781 + j-0.749084472656
            im_multiplicator=>-12273
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(748),
            data_im_in=>first_stage_im_out(748),
            product_re_out=>mul_re_out(748),
            product_im_out=>mul_im_out(748)
        );

    UMUL_749 : complex_multiplier
    generic map(
            re_multiplicator=>9960, --- 0.60791015625 + j-0.7939453125
            im_multiplicator=>-13008
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(749),
            data_im_in=>first_stage_im_out(749),
            product_re_out=>mul_re_out(749),
            product_im_out=>mul_im_out(749)
        );

    UMUL_750 : complex_multiplier
    generic map(
            re_multiplicator=>9018, --- 0.550415039062 + j-0.834838867188
            im_multiplicator=>-13678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(750),
            data_im_in=>first_stage_im_out(750),
            product_re_out=>mul_re_out(750),
            product_im_out=>mul_im_out(750)
        );

    UMUL_751 : complex_multiplier
    generic map(
            re_multiplicator=>8031, --- 0.490173339844 + j-0.87158203125
            im_multiplicator=>-14280
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(751),
            data_im_in=>first_stage_im_out(751),
            product_re_out=>mul_re_out(751),
            product_im_out=>mul_im_out(751)
        );

    UMUL_752 : complex_multiplier
    generic map(
            re_multiplicator=>7005, --- 0.427551269531 + j-0.903930664062
            im_multiplicator=>-14810
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(752),
            data_im_in=>first_stage_im_out(752),
            product_re_out=>mul_re_out(752),
            product_im_out=>mul_im_out(752)
        );

    UMUL_753 : complex_multiplier
    generic map(
            re_multiplicator=>5943, --- 0.362731933594 + j-0.931823730469
            im_multiplicator=>-15267
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(753),
            data_im_in=>first_stage_im_out(753),
            product_re_out=>mul_re_out(753),
            product_im_out=>mul_im_out(753)
        );

    UMUL_754 : complex_multiplier
    generic map(
            re_multiplicator=>4852, --- 0.296142578125 + j-0.955139160156
            im_multiplicator=>-15649
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(754),
            data_im_in=>first_stage_im_out(754),
            product_re_out=>mul_re_out(754),
            product_im_out=>mul_im_out(754)
        );

    UMUL_755 : complex_multiplier
    generic map(
            re_multiplicator=>3736, --- 0.22802734375 + j-0.9736328125
            im_multiplicator=>-15952
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(755),
            data_im_in=>first_stage_im_out(755),
            product_re_out=>mul_re_out(755),
            product_im_out=>mul_im_out(755)
        );

    UMUL_756 : complex_multiplier
    generic map(
            re_multiplicator=>2602, --- 0.158813476562 + j-0.987243652344
            im_multiplicator=>-16175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(756),
            data_im_in=>first_stage_im_out(756),
            product_re_out=>mul_re_out(756),
            product_im_out=>mul_im_out(756)
        );

    UMUL_757 : complex_multiplier
    generic map(
            re_multiplicator=>1455, --- 0.0888061523438 + j-0.996032714844
            im_multiplicator=>-16319
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(757),
            data_im_in=>first_stage_im_out(757),
            product_re_out=>mul_re_out(757),
            product_im_out=>mul_im_out(757)
        );

    UMUL_758 : complex_multiplier
    generic map(
            re_multiplicator=>301, --- 0.0183715820312 + j-0.999816894531
            im_multiplicator=>-16381
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(758),
            data_im_in=>first_stage_im_out(758),
            product_re_out=>mul_re_out(758),
            product_im_out=>mul_im_out(758)
        );

    UMUL_759 : complex_multiplier
    generic map(
            re_multiplicator=>-854, --- -0.0521240234375 + j-0.998596191406
            im_multiplicator=>-16361
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(759),
            data_im_in=>first_stage_im_out(759),
            product_re_out=>mul_re_out(759),
            product_im_out=>mul_im_out(759)
        );

    UMUL_760 : complex_multiplier
    generic map(
            re_multiplicator=>-2005, --- -0.122375488281 + j-0.992431640625
            im_multiplicator=>-16260
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(760),
            data_im_in=>first_stage_im_out(760),
            product_re_out=>mul_re_out(760),
            product_im_out=>mul_im_out(760)
        );

    UMUL_761 : complex_multiplier
    generic map(
            re_multiplicator=>-3147, --- -0.192077636719 + j-0.981323242188
            im_multiplicator=>-16078
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(761),
            data_im_in=>first_stage_im_out(761),
            product_re_out=>mul_re_out(761),
            product_im_out=>mul_im_out(761)
        );

    UMUL_762 : complex_multiplier
    generic map(
            re_multiplicator=>-4272, --- -0.2607421875 + j-0.965393066406
            im_multiplicator=>-15817
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(762),
            data_im_in=>first_stage_im_out(762),
            product_re_out=>mul_re_out(762),
            product_im_out=>mul_im_out(762)
        );

    UMUL_763 : complex_multiplier
    generic map(
            re_multiplicator=>-5377, --- -0.328186035156 + j-0.944580078125
            im_multiplicator=>-15476
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(763),
            data_im_in=>first_stage_im_out(763),
            product_re_out=>mul_re_out(763),
            product_im_out=>mul_im_out(763)
        );

    UMUL_764 : complex_multiplier
    generic map(
            re_multiplicator=>-6455, --- -0.393981933594 + j-0.919067382812
            im_multiplicator=>-15058
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(764),
            data_im_in=>first_stage_im_out(764),
            product_re_out=>mul_re_out(764),
            product_im_out=>mul_im_out(764)
        );

    UMUL_765 : complex_multiplier
    generic map(
            re_multiplicator=>-7500, --- -0.457763671875 + j-0.889038085938
            im_multiplicator=>-14566
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(765),
            data_im_in=>first_stage_im_out(765),
            product_re_out=>mul_re_out(765),
            product_im_out=>mul_im_out(765)
        );

    UMUL_766 : complex_multiplier
    generic map(
            re_multiplicator=>-8509, --- -0.519348144531 + j-0.854553222656
            im_multiplicator=>-14001
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(766),
            data_im_in=>first_stage_im_out(766),
            product_re_out=>mul_re_out(766),
            product_im_out=>mul_im_out(766)
        );

    UMUL_767 : complex_multiplier
    generic map(
            re_multiplicator=>-9475, --- -0.578308105469 + j-0.815795898438
            im_multiplicator=>-13366
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(767),
            data_im_in=>first_stage_im_out(767),
            product_re_out=>mul_re_out(767),
            product_im_out=>mul_im_out(767)
        );

    UDELAY_768_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(768),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(768)
        );
    UDELAY_768_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(768),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(768)
        );
    USHIFTER_768_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(768),
            data_out=>mul_re_out(768)
        );
    USHIFTER_768_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(768),
            data_out=>mul_im_out(768)
        );

    UMUL_769 : complex_multiplier
    generic map(
            re_multiplicator=>16339, --- 0.997253417969 + j-0.0735473632812
            im_multiplicator=>-1205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(769),
            data_im_in=>first_stage_im_out(769),
            product_re_out=>mul_re_out(769),
            product_im_out=>mul_im_out(769)
        );

    UMUL_770 : complex_multiplier
    generic map(
            re_multiplicator=>16206, --- 0.989135742188 + j-0.146728515625
            im_multiplicator=>-2404
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(770),
            data_im_in=>first_stage_im_out(770),
            product_re_out=>mul_re_out(770),
            product_im_out=>mul_im_out(770)
        );

    UMUL_771 : complex_multiplier
    generic map(
            re_multiplicator=>15985, --- 0.975646972656 + j-0.219055175781
            im_multiplicator=>-3589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(771),
            data_im_in=>first_stage_im_out(771),
            product_re_out=>mul_re_out(771),
            product_im_out=>mul_im_out(771)
        );

    UMUL_772 : complex_multiplier
    generic map(
            re_multiplicator=>15678, --- 0.956909179688 + j-0.290283203125
            im_multiplicator=>-4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(772),
            data_im_in=>first_stage_im_out(772),
            product_re_out=>mul_re_out(772),
            product_im_out=>mul_im_out(772)
        );

    UMUL_773 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(773),
            data_im_in=>first_stage_im_out(773),
            product_re_out=>mul_re_out(773),
            product_im_out=>mul_im_out(773)
        );

    UMUL_774 : complex_multiplier
    generic map(
            re_multiplicator=>14810, --- 0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(774),
            data_im_in=>first_stage_im_out(774),
            product_re_out=>mul_re_out(774),
            product_im_out=>mul_im_out(774)
        );

    UMUL_775 : complex_multiplier
    generic map(
            re_multiplicator=>14255, --- 0.870056152344 + j-0.492858886719
            im_multiplicator=>-8075
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(775),
            data_im_in=>first_stage_im_out(775),
            product_re_out=>mul_re_out(775),
            product_im_out=>mul_im_out(775)
        );

    UMUL_776 : complex_multiplier
    generic map(
            re_multiplicator=>13622, --- 0.831420898438 + j-0.555541992188
            im_multiplicator=>-9102
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(776),
            data_im_in=>first_stage_im_out(776),
            product_re_out=>mul_re_out(776),
            product_im_out=>mul_im_out(776)
        );

    UMUL_777 : complex_multiplier
    generic map(
            re_multiplicator=>12916, --- 0.788330078125 + j-0.615173339844
            im_multiplicator=>-10079
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(777),
            data_im_in=>first_stage_im_out(777),
            product_re_out=>mul_re_out(777),
            product_im_out=>mul_im_out(777)
        );

    UMUL_778 : complex_multiplier
    generic map(
            re_multiplicator=>12139, --- 0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(778),
            data_im_in=>first_stage_im_out(778),
            product_re_out=>mul_re_out(778),
            product_im_out=>mul_im_out(778)
        );

    UMUL_779 : complex_multiplier
    generic map(
            re_multiplicator=>11297, --- 0.689514160156 + j-0.724243164062
            im_multiplicator=>-11866
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(779),
            data_im_in=>first_stage_im_out(779),
            product_re_out=>mul_re_out(779),
            product_im_out=>mul_im_out(779)
        );

    UMUL_780 : complex_multiplier
    generic map(
            re_multiplicator=>10393, --- 0.634338378906 + j-0.773010253906
            im_multiplicator=>-12665
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(780),
            data_im_in=>first_stage_im_out(780),
            product_re_out=>mul_re_out(780),
            product_im_out=>mul_im_out(780)
        );

    UMUL_781 : complex_multiplier
    generic map(
            re_multiplicator=>9434, --- 0.575805664062 + j-0.817565917969
            im_multiplicator=>-13395
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(781),
            data_im_in=>first_stage_im_out(781),
            product_re_out=>mul_re_out(781),
            product_im_out=>mul_im_out(781)
        );

    UMUL_782 : complex_multiplier
    generic map(
            re_multiplicator=>8423, --- 0.514099121094 + j-0.857727050781
            im_multiplicator=>-14053
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(782),
            data_im_in=>first_stage_im_out(782),
            product_re_out=>mul_re_out(782),
            product_im_out=>mul_im_out(782)
        );

    UMUL_783 : complex_multiplier
    generic map(
            re_multiplicator=>7366, --- 0.449584960938 + j-0.893188476562
            im_multiplicator=>-14634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(783),
            data_im_in=>first_stage_im_out(783),
            product_re_out=>mul_re_out(783),
            product_im_out=>mul_im_out(783)
        );

    UMUL_784 : complex_multiplier
    generic map(
            re_multiplicator=>6269, --- 0.382629394531 + j-0.923828125
            im_multiplicator=>-15136
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(784),
            data_im_in=>first_stage_im_out(784),
            product_re_out=>mul_re_out(784),
            product_im_out=>mul_im_out(784)
        );

    UMUL_785 : complex_multiplier
    generic map(
            re_multiplicator=>5139, --- 0.313659667969 + j-0.949523925781
            im_multiplicator=>-15557
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(785),
            data_im_in=>first_stage_im_out(785),
            product_re_out=>mul_re_out(785),
            product_im_out=>mul_im_out(785)
        );

    UMUL_786 : complex_multiplier
    generic map(
            re_multiplicator=>3980, --- 0.242919921875 + j-0.969970703125
            im_multiplicator=>-15892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(786),
            data_im_in=>first_stage_im_out(786),
            product_re_out=>mul_re_out(786),
            product_im_out=>mul_im_out(786)
        );

    UMUL_787 : complex_multiplier
    generic map(
            re_multiplicator=>2801, --- 0.170959472656 + j-0.985229492188
            im_multiplicator=>-16142
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(787),
            data_im_in=>first_stage_im_out(787),
            product_re_out=>mul_re_out(787),
            product_im_out=>mul_im_out(787)
        );

    UMUL_788 : complex_multiplier
    generic map(
            re_multiplicator=>1605, --- 0.0979614257812 + j-0.995178222656
            im_multiplicator=>-16305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(788),
            data_im_in=>first_stage_im_out(788),
            product_re_out=>mul_re_out(788),
            product_im_out=>mul_im_out(788)
        );

    UMUL_789 : complex_multiplier
    generic map(
            re_multiplicator=>402, --- 0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(789),
            data_im_in=>first_stage_im_out(789),
            product_re_out=>mul_re_out(789),
            product_im_out=>mul_im_out(789)
        );

    UMUL_790 : complex_multiplier
    generic map(
            re_multiplicator=>-803, --- -0.0490112304688 + j-0.998779296875
            im_multiplicator=>-16364
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(790),
            data_im_in=>first_stage_im_out(790),
            product_re_out=>mul_re_out(790),
            product_im_out=>mul_im_out(790)
        );

    UMUL_791 : complex_multiplier
    generic map(
            re_multiplicator=>-2005, --- -0.122375488281 + j-0.992431640625
            im_multiplicator=>-16260
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(791),
            data_im_in=>first_stage_im_out(791),
            product_re_out=>mul_re_out(791),
            product_im_out=>mul_im_out(791)
        );

    UMUL_792 : complex_multiplier
    generic map(
            re_multiplicator=>-3196, --- -0.195068359375 + j-0.980773925781
            im_multiplicator=>-16069
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(792),
            data_im_in=>first_stage_im_out(792),
            product_re_out=>mul_re_out(792),
            product_im_out=>mul_im_out(792)
        );

    UMUL_793 : complex_multiplier
    generic map(
            re_multiplicator=>-4369, --- -0.266662597656 + j-0.963745117188
            im_multiplicator=>-15790
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(793),
            data_im_in=>first_stage_im_out(793),
            product_re_out=>mul_re_out(793),
            product_im_out=>mul_im_out(793)
        );

    UMUL_794 : complex_multiplier
    generic map(
            re_multiplicator=>-5519, --- -0.336853027344 + j-0.941528320312
            im_multiplicator=>-15426
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(794),
            data_im_in=>first_stage_im_out(794),
            product_re_out=>mul_re_out(794),
            product_im_out=>mul_im_out(794)
        );

    UMUL_795 : complex_multiplier
    generic map(
            re_multiplicator=>-6639, --- -0.405212402344 + j-0.914184570312
            im_multiplicator=>-14978
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(795),
            data_im_in=>first_stage_im_out(795),
            product_re_out=>mul_re_out(795),
            product_im_out=>mul_im_out(795)
        );

    UMUL_796 : complex_multiplier
    generic map(
            re_multiplicator=>-7723, --- -0.471374511719 + j-0.881896972656
            im_multiplicator=>-14449
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(796),
            data_im_in=>first_stage_im_out(796),
            product_re_out=>mul_re_out(796),
            product_im_out=>mul_im_out(796)
        );

    UMUL_797 : complex_multiplier
    generic map(
            re_multiplicator=>-8765, --- -0.534973144531 + j-0.844848632812
            im_multiplicator=>-13842
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(797),
            data_im_in=>first_stage_im_out(797),
            product_re_out=>mul_re_out(797),
            product_im_out=>mul_im_out(797)
        );

    UMUL_798 : complex_multiplier
    generic map(
            re_multiplicator=>-9759, --- -0.595642089844 + j-0.803161621094
            im_multiplicator=>-13159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(798),
            data_im_in=>first_stage_im_out(798),
            product_re_out=>mul_re_out(798),
            product_im_out=>mul_im_out(798)
        );

    UMUL_799 : complex_multiplier
    generic map(
            re_multiplicator=>-10701, --- -0.653137207031 + j-0.757202148438
            im_multiplicator=>-12406
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(799),
            data_im_in=>first_stage_im_out(799),
            product_re_out=>mul_re_out(799),
            product_im_out=>mul_im_out(799)
        );

    UDELAY_800_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(800),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(800)
        );
    UDELAY_800_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(800),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(800)
        );
    USHIFTER_800_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(800),
            data_out=>mul_re_out(800)
        );
    USHIFTER_800_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(800),
            data_out=>mul_im_out(800)
        );

    UMUL_801 : complex_multiplier
    generic map(
            re_multiplicator=>16335, --- 0.997009277344 + j-0.0765991210938
            im_multiplicator=>-1255
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(801),
            data_im_in=>first_stage_im_out(801),
            product_re_out=>mul_re_out(801),
            product_im_out=>mul_im_out(801)
        );

    UMUL_802 : complex_multiplier
    generic map(
            re_multiplicator=>16191, --- 0.988220214844 + j-0.152770996094
            im_multiplicator=>-2503
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(802),
            data_im_in=>first_stage_im_out(802),
            product_re_out=>mul_re_out(802),
            product_im_out=>mul_im_out(802)
        );

    UMUL_803 : complex_multiplier
    generic map(
            re_multiplicator=>15952, --- 0.9736328125 + j-0.22802734375
            im_multiplicator=>-3736
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(803),
            data_im_in=>first_stage_im_out(803),
            product_re_out=>mul_re_out(803),
            product_im_out=>mul_im_out(803)
        );

    UMUL_804 : complex_multiplier
    generic map(
            re_multiplicator=>15618, --- 0.953247070312 + j-0.302001953125
            im_multiplicator=>-4948
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(804),
            data_im_in=>first_stage_im_out(804),
            product_re_out=>mul_re_out(804),
            product_im_out=>mul_im_out(804)
        );

    UMUL_805 : complex_multiplier
    generic map(
            re_multiplicator=>15193, --- 0.927307128906 + j-0.374145507812
            im_multiplicator=>-6130
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(805),
            data_im_in=>first_stage_im_out(805),
            product_re_out=>mul_re_out(805),
            product_im_out=>mul_im_out(805)
        );

    UMUL_806 : complex_multiplier
    generic map(
            re_multiplicator=>14679, --- 0.895935058594 + j-0.444091796875
            im_multiplicator=>-7276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(806),
            data_im_in=>first_stage_im_out(806),
            product_re_out=>mul_re_out(806),
            product_im_out=>mul_im_out(806)
        );

    UMUL_807 : complex_multiplier
    generic map(
            re_multiplicator=>14078, --- 0.859252929688 + j-0.511413574219
            im_multiplicator=>-8379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(807),
            data_im_in=>first_stage_im_out(807),
            product_re_out=>mul_re_out(807),
            product_im_out=>mul_im_out(807)
        );

    UMUL_808 : complex_multiplier
    generic map(
            re_multiplicator=>13395, --- 0.817565917969 + j-0.575805664062
            im_multiplicator=>-9434
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(808),
            data_im_in=>first_stage_im_out(808),
            product_re_out=>mul_re_out(808),
            product_im_out=>mul_im_out(808)
        );

    UMUL_809 : complex_multiplier
    generic map(
            re_multiplicator=>12633, --- 0.771057128906 + j-0.63671875
            im_multiplicator=>-10432
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(809),
            data_im_in=>first_stage_im_out(809),
            product_re_out=>mul_re_out(809),
            product_im_out=>mul_im_out(809)
        );

    UMUL_810 : complex_multiplier
    generic map(
            re_multiplicator=>11796, --- 0.719970703125 + j-0.693969726562
            im_multiplicator=>-11370
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(810),
            data_im_in=>first_stage_im_out(810),
            product_re_out=>mul_re_out(810),
            product_im_out=>mul_im_out(810)
        );

    UMUL_811 : complex_multiplier
    generic map(
            re_multiplicator=>10890, --- 0.664672851562 + j-0.7470703125
            im_multiplicator=>-12240
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(811),
            data_im_in=>first_stage_im_out(811),
            product_re_out=>mul_re_out(811),
            product_im_out=>mul_im_out(811)
        );

    UMUL_812 : complex_multiplier
    generic map(
            re_multiplicator=>9920, --- 0.60546875 + j-0.795776367188
            im_multiplicator=>-13038
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(812),
            data_im_in=>first_stage_im_out(812),
            product_re_out=>mul_re_out(812),
            product_im_out=>mul_im_out(812)
        );

    UMUL_813 : complex_multiplier
    generic map(
            re_multiplicator=>8892, --- 0.542724609375 + j-0.83984375
            im_multiplicator=>-13760
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(813),
            data_im_in=>first_stage_im_out(813),
            product_re_out=>mul_re_out(813),
            product_im_out=>mul_im_out(813)
        );

    UMUL_814 : complex_multiplier
    generic map(
            re_multiplicator=>7811, --- 0.476745605469 + j-0.878967285156
            im_multiplicator=>-14401
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(814),
            data_im_in=>first_stage_im_out(814),
            product_re_out=>mul_re_out(814),
            product_im_out=>mul_im_out(814)
        );

    UMUL_815 : complex_multiplier
    generic map(
            re_multiplicator=>6685, --- 0.408020019531 + j-0.912902832031
            im_multiplicator=>-14957
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(815),
            data_im_in=>first_stage_im_out(815),
            product_re_out=>mul_re_out(815),
            product_im_out=>mul_im_out(815)
        );

    UMUL_816 : complex_multiplier
    generic map(
            re_multiplicator=>5519, --- 0.336853027344 + j-0.941528320312
            im_multiplicator=>-15426
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(816),
            data_im_in=>first_stage_im_out(816),
            product_re_out=>mul_re_out(816),
            product_im_out=>mul_im_out(816)
        );

    UMUL_817 : complex_multiplier
    generic map(
            re_multiplicator=>4321, --- 0.263732910156 + j-0.964538574219
            im_multiplicator=>-15803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(817),
            data_im_in=>first_stage_im_out(817),
            product_re_out=>mul_re_out(817),
            product_im_out=>mul_im_out(817)
        );

    UMUL_818 : complex_multiplier
    generic map(
            re_multiplicator=>3097, --- 0.189025878906 + j-0.98193359375
            im_multiplicator=>-16088
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(818),
            data_im_in=>first_stage_im_out(818),
            product_re_out=>mul_re_out(818),
            product_im_out=>mul_im_out(818)
        );

    UMUL_819 : complex_multiplier
    generic map(
            re_multiplicator=>1855, --- 0.113220214844 + j-0.993530273438
            im_multiplicator=>-16278
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(819),
            data_im_in=>first_stage_im_out(819),
            product_re_out=>mul_re_out(819),
            product_im_out=>mul_im_out(819)
        );

    UMUL_820 : complex_multiplier
    generic map(
            re_multiplicator=>603, --- 0.0368041992188 + j-0.999267578125
            im_multiplicator=>-16372
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(820),
            data_im_in=>first_stage_im_out(820),
            product_re_out=>mul_re_out(820),
            product_im_out=>mul_im_out(820)
        );

    UMUL_821 : complex_multiplier
    generic map(
            re_multiplicator=>-653, --- -0.0398559570312 + j-0.999145507812
            im_multiplicator=>-16370
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(821),
            data_im_in=>first_stage_im_out(821),
            product_re_out=>mul_re_out(821),
            product_im_out=>mul_im_out(821)
        );

    UMUL_822 : complex_multiplier
    generic map(
            re_multiplicator=>-1905, --- -0.116271972656 + j-0.9931640625
            im_multiplicator=>-16272
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(822),
            data_im_in=>first_stage_im_out(822),
            product_re_out=>mul_re_out(822),
            product_im_out=>mul_im_out(822)
        );

    UMUL_823 : complex_multiplier
    generic map(
            re_multiplicator=>-3147, --- -0.192077636719 + j-0.981323242188
            im_multiplicator=>-16078
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(823),
            data_im_in=>first_stage_im_out(823),
            product_re_out=>mul_re_out(823),
            product_im_out=>mul_im_out(823)
        );

    UMUL_824 : complex_multiplier
    generic map(
            re_multiplicator=>-4369, --- -0.266662597656 + j-0.963745117188
            im_multiplicator=>-15790
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(824),
            data_im_in=>first_stage_im_out(824),
            product_re_out=>mul_re_out(824),
            product_im_out=>mul_im_out(824)
        );

    UMUL_825 : complex_multiplier
    generic map(
            re_multiplicator=>-5566, --- -0.339721679688 + j-0.940490722656
            im_multiplicator=>-15409
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(825),
            data_im_in=>first_stage_im_out(825),
            product_re_out=>mul_re_out(825),
            product_im_out=>mul_im_out(825)
        );

    UMUL_826 : complex_multiplier
    generic map(
            re_multiplicator=>-6731, --- -0.410827636719 + j-0.911682128906
            im_multiplicator=>-14937
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(826),
            data_im_in=>first_stage_im_out(826),
            product_re_out=>mul_re_out(826),
            product_im_out=>mul_im_out(826)
        );

    UMUL_827 : complex_multiplier
    generic map(
            re_multiplicator=>-7856, --- -0.4794921875 + j-0.877502441406
            im_multiplicator=>-14377
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(827),
            data_im_in=>first_stage_im_out(827),
            product_re_out=>mul_re_out(827),
            product_im_out=>mul_im_out(827)
        );

    UMUL_828 : complex_multiplier
    generic map(
            re_multiplicator=>-8934, --- -0.545288085938 + j-0.838195800781
            im_multiplicator=>-13733
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(828),
            data_im_in=>first_stage_im_out(828),
            product_re_out=>mul_re_out(828),
            product_im_out=>mul_im_out(828)
        );

    UMUL_829 : complex_multiplier
    generic map(
            re_multiplicator=>-9960, --- -0.60791015625 + j-0.7939453125
            im_multiplicator=>-13008
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(829),
            data_im_in=>first_stage_im_out(829),
            product_re_out=>mul_re_out(829),
            product_im_out=>mul_im_out(829)
        );

    UMUL_830 : complex_multiplier
    generic map(
            re_multiplicator=>-10928, --- -0.6669921875 + j-0.745056152344
            im_multiplicator=>-12207
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(830),
            data_im_in=>first_stage_im_out(830),
            product_re_out=>mul_re_out(830),
            product_im_out=>mul_im_out(830)
        );

    UMUL_831 : complex_multiplier
    generic map(
            re_multiplicator=>-11831, --- -0.722106933594 + j-0.691711425781
            im_multiplicator=>-11333
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(831),
            data_im_in=>first_stage_im_out(831),
            product_re_out=>mul_re_out(831),
            product_im_out=>mul_im_out(831)
        );

    UDELAY_832_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(832),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(832)
        );
    UDELAY_832_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(832),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(832)
        );
    USHIFTER_832_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(832),
            data_out=>mul_re_out(832)
        );
    USHIFTER_832_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(832),
            data_out=>mul_im_out(832)
        );

    UMUL_833 : complex_multiplier
    generic map(
            re_multiplicator=>16331, --- 0.996765136719 + j-0.0796508789062
            im_multiplicator=>-1305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(833),
            data_im_in=>first_stage_im_out(833),
            product_re_out=>mul_re_out(833),
            product_im_out=>mul_im_out(833)
        );

    UMUL_834 : complex_multiplier
    generic map(
            re_multiplicator=>16175, --- 0.987243652344 + j-0.158813476562
            im_multiplicator=>-2602
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(834),
            data_im_in=>first_stage_im_out(834),
            product_re_out=>mul_re_out(834),
            product_im_out=>mul_im_out(834)
        );

    UMUL_835 : complex_multiplier
    generic map(
            re_multiplicator=>15917, --- 0.971496582031 + j-0.236999511719
            im_multiplicator=>-3883
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(835),
            data_im_in=>first_stage_im_out(835),
            product_re_out=>mul_re_out(835),
            product_im_out=>mul_im_out(835)
        );

    UMUL_836 : complex_multiplier
    generic map(
            re_multiplicator=>15557, --- 0.949523925781 + j-0.313659667969
            im_multiplicator=>-5139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(836),
            data_im_in=>first_stage_im_out(836),
            product_re_out=>mul_re_out(836),
            product_im_out=>mul_im_out(836)
        );

    UMUL_837 : complex_multiplier
    generic map(
            re_multiplicator=>15098, --- 0.921508789062 + j-0.388305664062
            im_multiplicator=>-6362
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(837),
            data_im_in=>first_stage_im_out(837),
            product_re_out=>mul_re_out(837),
            product_im_out=>mul_im_out(837)
        );

    UMUL_838 : complex_multiplier
    generic map(
            re_multiplicator=>14543, --- 0.887634277344 + j-0.460510253906
            im_multiplicator=>-7545
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(838),
            data_im_in=>first_stage_im_out(838),
            product_re_out=>mul_re_out(838),
            product_im_out=>mul_im_out(838)
        );

    UMUL_839 : complex_multiplier
    generic map(
            re_multiplicator=>13895, --- 0.848083496094 + j-0.52978515625
            im_multiplicator=>-8680
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(839),
            data_im_in=>first_stage_im_out(839),
            product_re_out=>mul_re_out(839),
            product_im_out=>mul_im_out(839)
        );

    UMUL_840 : complex_multiplier
    generic map(
            re_multiplicator=>13159, --- 0.803161621094 + j-0.595642089844
            im_multiplicator=>-9759
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(840),
            data_im_in=>first_stage_im_out(840),
            product_re_out=>mul_re_out(840),
            product_im_out=>mul_im_out(840)
        );

    UMUL_841 : complex_multiplier
    generic map(
            re_multiplicator=>12340, --- 0.753173828125 + j-0.657775878906
            im_multiplicator=>-10777
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(841),
            data_im_in=>first_stage_im_out(841),
            product_re_out=>mul_re_out(841),
            product_im_out=>mul_im_out(841)
        );

    UMUL_842 : complex_multiplier
    generic map(
            re_multiplicator=>11442, --- 0.698364257812 + j-0.715698242188
            im_multiplicator=>-11726
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(842),
            data_im_in=>first_stage_im_out(842),
            product_re_out=>mul_re_out(842),
            product_im_out=>mul_im_out(842)
        );

    UMUL_843 : complex_multiplier
    generic map(
            re_multiplicator=>10471, --- 0.639099121094 + j-0.76904296875
            im_multiplicator=>-12600
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(843),
            data_im_in=>first_stage_im_out(843),
            product_re_out=>mul_re_out(843),
            product_im_out=>mul_im_out(843)
        );

    UMUL_844 : complex_multiplier
    generic map(
            re_multiplicator=>9434, --- 0.575805664062 + j-0.817565917969
            im_multiplicator=>-13395
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(844),
            data_im_in=>first_stage_im_out(844),
            product_re_out=>mul_re_out(844),
            product_im_out=>mul_im_out(844)
        );

    UMUL_845 : complex_multiplier
    generic map(
            re_multiplicator=>8336, --- 0.5087890625 + j-0.86083984375
            im_multiplicator=>-14104
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(845),
            data_im_in=>first_stage_im_out(845),
            product_re_out=>mul_re_out(845),
            product_im_out=>mul_im_out(845)
        );

    UMUL_846 : complex_multiplier
    generic map(
            re_multiplicator=>7186, --- 0.438598632812 + j-0.898620605469
            im_multiplicator=>-14723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(846),
            data_im_in=>first_stage_im_out(846),
            product_re_out=>mul_re_out(846),
            product_im_out=>mul_im_out(846)
        );

    UMUL_847 : complex_multiplier
    generic map(
            re_multiplicator=>5990, --- 0.365600585938 + j-0.930725097656
            im_multiplicator=>-15249
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(847),
            data_im_in=>first_stage_im_out(847),
            product_re_out=>mul_re_out(847),
            product_im_out=>mul_im_out(847)
        );

    UMUL_848 : complex_multiplier
    generic map(
            re_multiplicator=>4756, --- 0.290283203125 + j-0.956909179688
            im_multiplicator=>-15678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(848),
            data_im_in=>first_stage_im_out(848),
            product_re_out=>mul_re_out(848),
            product_im_out=>mul_im_out(848)
        );

    UMUL_849 : complex_multiplier
    generic map(
            re_multiplicator=>3491, --- 0.213073730469 + j-0.976989746094
            im_multiplicator=>-16007
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(849),
            data_im_in=>first_stage_im_out(849),
            product_re_out=>mul_re_out(849),
            product_im_out=>mul_im_out(849)
        );

    UMUL_850 : complex_multiplier
    generic map(
            re_multiplicator=>2204, --- 0.134521484375 + j-0.990844726562
            im_multiplicator=>-16234
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(850),
            data_im_in=>first_stage_im_out(850),
            product_re_out=>mul_re_out(850),
            product_im_out=>mul_im_out(850)
        );

    UMUL_851 : complex_multiplier
    generic map(
            re_multiplicator=>904, --- 0.05517578125 + j-0.998474121094
            im_multiplicator=>-16359
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(851),
            data_im_in=>first_stage_im_out(851),
            product_re_out=>mul_re_out(851),
            product_im_out=>mul_im_out(851)
        );

    UMUL_852 : complex_multiplier
    generic map(
            re_multiplicator=>-402, --- -0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(852),
            data_im_in=>first_stage_im_out(852),
            product_re_out=>mul_re_out(852),
            product_im_out=>mul_im_out(852)
        );

    UMUL_853 : complex_multiplier
    generic map(
            re_multiplicator=>-1705, --- -0.104064941406 + j-0.994506835938
            im_multiplicator=>-16294
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(853),
            data_im_in=>first_stage_im_out(853),
            product_re_out=>mul_re_out(853),
            product_im_out=>mul_im_out(853)
        );

    UMUL_854 : complex_multiplier
    generic map(
            re_multiplicator=>-2998, --- -0.182983398438 + j-0.983093261719
            im_multiplicator=>-16107
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(854),
            data_im_in=>first_stage_im_out(854),
            product_re_out=>mul_re_out(854),
            product_im_out=>mul_im_out(854)
        );

    UMUL_855 : complex_multiplier
    generic map(
            re_multiplicator=>-4272, --- -0.2607421875 + j-0.965393066406
            im_multiplicator=>-15817
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(855),
            data_im_in=>first_stage_im_out(855),
            product_re_out=>mul_re_out(855),
            product_im_out=>mul_im_out(855)
        );

    UMUL_856 : complex_multiplier
    generic map(
            re_multiplicator=>-5519, --- -0.336853027344 + j-0.941528320312
            im_multiplicator=>-15426
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(856),
            data_im_in=>first_stage_im_out(856),
            product_re_out=>mul_re_out(856),
            product_im_out=>mul_im_out(856)
        );

    UMUL_857 : complex_multiplier
    generic map(
            re_multiplicator=>-6731, --- -0.410827636719 + j-0.911682128906
            im_multiplicator=>-14937
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(857),
            data_im_in=>first_stage_im_out(857),
            product_re_out=>mul_re_out(857),
            product_im_out=>mul_im_out(857)
        );

    UMUL_858 : complex_multiplier
    generic map(
            re_multiplicator=>-7900, --- -0.482177734375 + j-0.876037597656
            im_multiplicator=>-14353
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(858),
            data_im_in=>first_stage_im_out(858),
            product_re_out=>mul_re_out(858),
            product_im_out=>mul_im_out(858)
        );

    UMUL_859 : complex_multiplier
    generic map(
            re_multiplicator=>-9018, --- -0.550415039062 + j-0.834838867188
            im_multiplicator=>-13678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(859),
            data_im_in=>first_stage_im_out(859),
            product_re_out=>mul_re_out(859),
            product_im_out=>mul_im_out(859)
        );

    UMUL_860 : complex_multiplier
    generic map(
            re_multiplicator=>-10079, --- -0.615173339844 + j-0.788330078125
            im_multiplicator=>-12916
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(860),
            data_im_in=>first_stage_im_out(860),
            product_re_out=>mul_re_out(860),
            product_im_out=>mul_im_out(860)
        );

    UMUL_861 : complex_multiplier
    generic map(
            re_multiplicator=>-11077, --- -0.676086425781 + j-0.73681640625
            im_multiplicator=>-12072
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(861),
            data_im_in=>first_stage_im_out(861),
            product_re_out=>mul_re_out(861),
            product_im_out=>mul_im_out(861)
        );

    UMUL_862 : complex_multiplier
    generic map(
            re_multiplicator=>-12003, --- -0.732604980469 + j-0.680541992188
            im_multiplicator=>-11150
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(862),
            data_im_in=>first_stage_im_out(862),
            product_re_out=>mul_re_out(862),
            product_im_out=>mul_im_out(862)
        );

    UMUL_863 : complex_multiplier
    generic map(
            re_multiplicator=>-12854, --- -0.784545898438 + j-0.620056152344
            im_multiplicator=>-10159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(863),
            data_im_in=>first_stage_im_out(863),
            product_re_out=>mul_re_out(863),
            product_im_out=>mul_im_out(863)
        );

    UDELAY_864_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(864),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(864)
        );
    UDELAY_864_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(864),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(864)
        );
    USHIFTER_864_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(864),
            data_out=>mul_re_out(864)
        );
    USHIFTER_864_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(864),
            data_out=>mul_im_out(864)
        );

    UMUL_865 : complex_multiplier
    generic map(
            re_multiplicator=>16327, --- 0.996520996094 + j-0.0827026367188
            im_multiplicator=>-1355
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(865),
            data_im_in=>first_stage_im_out(865),
            product_re_out=>mul_re_out(865),
            product_im_out=>mul_im_out(865)
        );

    UMUL_866 : complex_multiplier
    generic map(
            re_multiplicator=>16159, --- 0.986267089844 + j-0.164855957031
            im_multiplicator=>-2701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(866),
            data_im_in=>first_stage_im_out(866),
            product_re_out=>mul_re_out(866),
            product_im_out=>mul_im_out(866)
        );

    UMUL_867 : complex_multiplier
    generic map(
            re_multiplicator=>15880, --- 0.96923828125 + j-0.245910644531
            im_multiplicator=>-4029
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(867),
            data_im_in=>first_stage_im_out(867),
            product_re_out=>mul_re_out(867),
            product_im_out=>mul_im_out(867)
        );

    UMUL_868 : complex_multiplier
    generic map(
            re_multiplicator=>15492, --- 0.945556640625 + j-0.325256347656
            im_multiplicator=>-5329
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(868),
            data_im_in=>first_stage_im_out(868),
            product_re_out=>mul_re_out(868),
            product_im_out=>mul_im_out(868)
        );

    UMUL_869 : complex_multiplier
    generic map(
            re_multiplicator=>14998, --- 0.915405273438 + j-0.402404785156
            im_multiplicator=>-6593
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(869),
            data_im_in=>first_stage_im_out(869),
            product_re_out=>mul_re_out(869),
            product_im_out=>mul_im_out(869)
        );

    UMUL_870 : complex_multiplier
    generic map(
            re_multiplicator=>14401, --- 0.878967285156 + j-0.476745605469
            im_multiplicator=>-7811
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(870),
            data_im_in=>first_stage_im_out(870),
            product_re_out=>mul_re_out(870),
            product_im_out=>mul_im_out(870)
        );

    UMUL_871 : complex_multiplier
    generic map(
            re_multiplicator=>13705, --- 0.836486816406 + j-0.5478515625
            im_multiplicator=>-8976
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(871),
            data_im_in=>first_stage_im_out(871),
            product_re_out=>mul_re_out(871),
            product_im_out=>mul_im_out(871)
        );

    UMUL_872 : complex_multiplier
    generic map(
            re_multiplicator=>12916, --- 0.788330078125 + j-0.615173339844
            im_multiplicator=>-10079
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(872),
            data_im_in=>first_stage_im_out(872),
            product_re_out=>mul_re_out(872),
            product_im_out=>mul_im_out(872)
        );

    UMUL_873 : complex_multiplier
    generic map(
            re_multiplicator=>12037, --- 0.734680175781 + j-0.678344726562
            im_multiplicator=>-11114
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(873),
            data_im_in=>first_stage_im_out(873),
            product_re_out=>mul_re_out(873),
            product_im_out=>mul_im_out(873)
        );

    UMUL_874 : complex_multiplier
    generic map(
            re_multiplicator=>11077, --- 0.676086425781 + j-0.73681640625
            im_multiplicator=>-12072
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(874),
            data_im_in=>first_stage_im_out(874),
            product_re_out=>mul_re_out(874),
            product_im_out=>mul_im_out(874)
        );

    UMUL_875 : complex_multiplier
    generic map(
            re_multiplicator=>10040, --- 0.61279296875 + j-0.790222167969
            im_multiplicator=>-12947
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(875),
            data_im_in=>first_stage_im_out(875),
            product_re_out=>mul_re_out(875),
            product_im_out=>mul_im_out(875)
        );

    UMUL_876 : complex_multiplier
    generic map(
            re_multiplicator=>8934, --- 0.545288085938 + j-0.838195800781
            im_multiplicator=>-13733
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(876),
            data_im_in=>first_stage_im_out(876),
            product_re_out=>mul_re_out(876),
            product_im_out=>mul_im_out(876)
        );

    UMUL_877 : complex_multiplier
    generic map(
            re_multiplicator=>7767, --- 0.474060058594 + j-0.880432128906
            im_multiplicator=>-14425
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(877),
            data_im_in=>first_stage_im_out(877),
            product_re_out=>mul_re_out(877),
            product_im_out=>mul_im_out(877)
        );

    UMUL_878 : complex_multiplier
    generic map(
            re_multiplicator=>6547, --- 0.399597167969 + j-0.916625976562
            im_multiplicator=>-15018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(878),
            data_im_in=>first_stage_im_out(878),
            product_re_out=>mul_re_out(878),
            product_im_out=>mul_im_out(878)
        );

    UMUL_879 : complex_multiplier
    generic map(
            re_multiplicator=>5282, --- 0.322387695312 + j-0.946594238281
            im_multiplicator=>-15509
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(879),
            data_im_in=>first_stage_im_out(879),
            product_re_out=>mul_re_out(879),
            product_im_out=>mul_im_out(879)
        );

    UMUL_880 : complex_multiplier
    generic map(
            re_multiplicator=>3980, --- 0.242919921875 + j-0.969970703125
            im_multiplicator=>-15892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(880),
            data_im_in=>first_stage_im_out(880),
            product_re_out=>mul_re_out(880),
            product_im_out=>mul_im_out(880)
        );

    UMUL_881 : complex_multiplier
    generic map(
            re_multiplicator=>2652, --- 0.161865234375 + j-0.986755371094
            im_multiplicator=>-16167
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(881),
            data_im_in=>first_stage_im_out(881),
            product_re_out=>mul_re_out(881),
            product_im_out=>mul_im_out(881)
        );

    UMUL_882 : complex_multiplier
    generic map(
            re_multiplicator=>1305, --- 0.0796508789062 + j-0.996765136719
            im_multiplicator=>-16331
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(882),
            data_im_in=>first_stage_im_out(882),
            product_re_out=>mul_re_out(882),
            product_im_out=>mul_im_out(882)
        );

    UMUL_883 : complex_multiplier
    generic map(
            re_multiplicator=>-50, --- -0.0030517578125 + j-0.999938964844
            im_multiplicator=>-16383
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(883),
            data_im_in=>first_stage_im_out(883),
            product_re_out=>mul_re_out(883),
            product_im_out=>mul_im_out(883)
        );

    UMUL_884 : complex_multiplier
    generic map(
            re_multiplicator=>-1405, --- -0.0857543945312 + j-0.996276855469
            im_multiplicator=>-16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(884),
            data_im_in=>first_stage_im_out(884),
            product_re_out=>mul_re_out(884),
            product_im_out=>mul_im_out(884)
        );

    UMUL_885 : complex_multiplier
    generic map(
            re_multiplicator=>-2751, --- -0.167907714844 + j-0.985778808594
            im_multiplicator=>-16151
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(885),
            data_im_in=>first_stage_im_out(885),
            product_re_out=>mul_re_out(885),
            product_im_out=>mul_im_out(885)
        );

    UMUL_886 : complex_multiplier
    generic map(
            re_multiplicator=>-4078, --- -0.248901367188 + j-0.968505859375
            im_multiplicator=>-15868
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(886),
            data_im_in=>first_stage_im_out(886),
            product_re_out=>mul_re_out(886),
            product_im_out=>mul_im_out(886)
        );

    UMUL_887 : complex_multiplier
    generic map(
            re_multiplicator=>-5377, --- -0.328186035156 + j-0.944580078125
            im_multiplicator=>-15476
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(887),
            data_im_in=>first_stage_im_out(887),
            product_re_out=>mul_re_out(887),
            product_im_out=>mul_im_out(887)
        );

    UMUL_888 : complex_multiplier
    generic map(
            re_multiplicator=>-6639, --- -0.405212402344 + j-0.914184570312
            im_multiplicator=>-14978
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(888),
            data_im_in=>first_stage_im_out(888),
            product_re_out=>mul_re_out(888),
            product_im_out=>mul_im_out(888)
        );

    UMUL_889 : complex_multiplier
    generic map(
            re_multiplicator=>-7856, --- -0.4794921875 + j-0.877502441406
            im_multiplicator=>-14377
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(889),
            data_im_in=>first_stage_im_out(889),
            product_re_out=>mul_re_out(889),
            product_im_out=>mul_im_out(889)
        );

    UMUL_890 : complex_multiplier
    generic map(
            re_multiplicator=>-9018, --- -0.550415039062 + j-0.834838867188
            im_multiplicator=>-13678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(890),
            data_im_in=>first_stage_im_out(890),
            product_re_out=>mul_re_out(890),
            product_im_out=>mul_im_out(890)
        );

    UMUL_891 : complex_multiplier
    generic map(
            re_multiplicator=>-10119, --- -0.617614746094 + j-0.786437988281
            im_multiplicator=>-12885
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(891),
            data_im_in=>first_stage_im_out(891),
            product_re_out=>mul_re_out(891),
            product_im_out=>mul_im_out(891)
        );

    UMUL_892 : complex_multiplier
    generic map(
            re_multiplicator=>-11150, --- -0.680541992188 + j-0.732604980469
            im_multiplicator=>-12003
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(892),
            data_im_in=>first_stage_im_out(892),
            product_re_out=>mul_re_out(892),
            product_im_out=>mul_im_out(892)
        );

    UMUL_893 : complex_multiplier
    generic map(
            re_multiplicator=>-12105, --- -0.738830566406 + j-0.673828125
            im_multiplicator=>-11040
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(893),
            data_im_in=>first_stage_im_out(893),
            product_re_out=>mul_re_out(893),
            product_im_out=>mul_im_out(893)
        );

    UMUL_894 : complex_multiplier
    generic map(
            re_multiplicator=>-12977, --- -0.792053222656 + j-0.6103515625
            im_multiplicator=>-10000
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(894),
            data_im_in=>first_stage_im_out(894),
            product_re_out=>mul_re_out(894),
            product_im_out=>mul_im_out(894)
        );

    UMUL_895 : complex_multiplier
    generic map(
            re_multiplicator=>-13760, --- -0.83984375 + j-0.542724609375
            im_multiplicator=>-8892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(895),
            data_im_in=>first_stage_im_out(895),
            product_re_out=>mul_re_out(895),
            product_im_out=>mul_im_out(895)
        );

    UDELAY_896_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(896),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(896)
        );
    UDELAY_896_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(896),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(896)
        );
    USHIFTER_896_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(896),
            data_out=>mul_re_out(896)
        );
    USHIFTER_896_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(896),
            data_out=>mul_im_out(896)
        );

    UMUL_897 : complex_multiplier
    generic map(
            re_multiplicator=>16323, --- 0.996276855469 + j-0.0857543945312
            im_multiplicator=>-1405
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(897),
            data_im_in=>first_stage_im_out(897),
            product_re_out=>mul_re_out(897),
            product_im_out=>mul_im_out(897)
        );

    UMUL_898 : complex_multiplier
    generic map(
            re_multiplicator=>16142, --- 0.985229492188 + j-0.170959472656
            im_multiplicator=>-2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(898),
            data_im_in=>first_stage_im_out(898),
            product_re_out=>mul_re_out(898),
            product_im_out=>mul_im_out(898)
        );

    UMUL_899 : complex_multiplier
    generic map(
            re_multiplicator=>15842, --- 0.966918945312 + j-0.254821777344
            im_multiplicator=>-4175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(899),
            data_im_in=>first_stage_im_out(899),
            product_re_out=>mul_re_out(899),
            product_im_out=>mul_im_out(899)
        );

    UMUL_900 : complex_multiplier
    generic map(
            re_multiplicator=>15426, --- 0.941528320312 + j-0.336853027344
            im_multiplicator=>-5519
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(900),
            data_im_in=>first_stage_im_out(900),
            product_re_out=>mul_re_out(900),
            product_im_out=>mul_im_out(900)
        );

    UMUL_901 : complex_multiplier
    generic map(
            re_multiplicator=>14895, --- 0.909118652344 + j-0.416381835938
            im_multiplicator=>-6822
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(901),
            data_im_in=>first_stage_im_out(901),
            product_re_out=>mul_re_out(901),
            product_im_out=>mul_im_out(901)
        );

    UMUL_902 : complex_multiplier
    generic map(
            re_multiplicator=>14255, --- 0.870056152344 + j-0.492858886719
            im_multiplicator=>-8075
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(902),
            data_im_in=>first_stage_im_out(902),
            product_re_out=>mul_re_out(902),
            product_im_out=>mul_im_out(902)
        );

    UMUL_903 : complex_multiplier
    generic map(
            re_multiplicator=>13510, --- 0.824584960938 + j-0.565673828125
            im_multiplicator=>-9268
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(903),
            data_im_in=>first_stage_im_out(903),
            product_re_out=>mul_re_out(903),
            product_im_out=>mul_im_out(903)
        );

    UMUL_904 : complex_multiplier
    generic map(
            re_multiplicator=>12665, --- 0.773010253906 + j-0.634338378906
            im_multiplicator=>-10393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(904),
            data_im_in=>first_stage_im_out(904),
            product_re_out=>mul_re_out(904),
            product_im_out=>mul_im_out(904)
        );

    UMUL_905 : complex_multiplier
    generic map(
            re_multiplicator=>11726, --- 0.715698242188 + j-0.698364257812
            im_multiplicator=>-11442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(905),
            data_im_in=>first_stage_im_out(905),
            product_re_out=>mul_re_out(905),
            product_im_out=>mul_im_out(905)
        );

    UMUL_906 : complex_multiplier
    generic map(
            re_multiplicator=>10701, --- 0.653137207031 + j-0.757202148438
            im_multiplicator=>-12406
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(906),
            data_im_in=>first_stage_im_out(906),
            product_re_out=>mul_re_out(906),
            product_im_out=>mul_im_out(906)
        );

    UMUL_907 : complex_multiplier
    generic map(
            re_multiplicator=>9597, --- 0.585754394531 + j-0.810424804688
            im_multiplicator=>-13278
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(907),
            data_im_in=>first_stage_im_out(907),
            product_re_out=>mul_re_out(907),
            product_im_out=>mul_im_out(907)
        );

    UMUL_908 : complex_multiplier
    generic map(
            re_multiplicator=>8423, --- 0.514099121094 + j-0.857727050781
            im_multiplicator=>-14053
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(908),
            data_im_in=>first_stage_im_out(908),
            product_re_out=>mul_re_out(908),
            product_im_out=>mul_im_out(908)
        );

    UMUL_909 : complex_multiplier
    generic map(
            re_multiplicator=>7186, --- 0.438598632812 + j-0.898620605469
            im_multiplicator=>-14723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(909),
            data_im_in=>first_stage_im_out(909),
            product_re_out=>mul_re_out(909),
            product_im_out=>mul_im_out(909)
        );

    UMUL_910 : complex_multiplier
    generic map(
            re_multiplicator=>5896, --- 0.35986328125 + j-0.932983398438
            im_multiplicator=>-15286
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(910),
            data_im_in=>first_stage_im_out(910),
            product_re_out=>mul_re_out(910),
            product_im_out=>mul_im_out(910)
        );

    UMUL_911 : complex_multiplier
    generic map(
            re_multiplicator=>4563, --- 0.278503417969 + j-0.960388183594
            im_multiplicator=>-15735
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(911),
            data_im_in=>first_stage_im_out(911),
            product_re_out=>mul_re_out(911),
            product_im_out=>mul_im_out(911)
        );

    UMUL_912 : complex_multiplier
    generic map(
            re_multiplicator=>3196, --- 0.195068359375 + j-0.980773925781
            im_multiplicator=>-16069
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(912),
            data_im_in=>first_stage_im_out(912),
            product_re_out=>mul_re_out(912),
            product_im_out=>mul_im_out(912)
        );

    UMUL_913 : complex_multiplier
    generic map(
            re_multiplicator=>1805, --- 0.110168457031 + j-0.993896484375
            im_multiplicator=>-16284
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(913),
            data_im_in=>first_stage_im_out(913),
            product_re_out=>mul_re_out(913),
            product_im_out=>mul_im_out(913)
        );

    UMUL_914 : complex_multiplier
    generic map(
            re_multiplicator=>402, --- 0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(914),
            data_im_in=>first_stage_im_out(914),
            product_re_out=>mul_re_out(914),
            product_im_out=>mul_im_out(914)
        );

    UMUL_915 : complex_multiplier
    generic map(
            re_multiplicator=>-1004, --- -0.061279296875 + j-0.998107910156
            im_multiplicator=>-16353
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(915),
            data_im_in=>first_stage_im_out(915),
            product_re_out=>mul_re_out(915),
            product_im_out=>mul_im_out(915)
        );

    UMUL_916 : complex_multiplier
    generic map(
            re_multiplicator=>-2404, --- -0.146728515625 + j-0.989135742188
            im_multiplicator=>-16206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(916),
            data_im_in=>first_stage_im_out(916),
            product_re_out=>mul_re_out(916),
            product_im_out=>mul_im_out(916)
        );

    UMUL_917 : complex_multiplier
    generic map(
            re_multiplicator=>-3785, --- -0.231018066406 + j-0.972900390625
            im_multiplicator=>-15940
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(917),
            data_im_in=>first_stage_im_out(917),
            product_re_out=>mul_re_out(917),
            product_im_out=>mul_im_out(917)
        );

    UMUL_918 : complex_multiplier
    generic map(
            re_multiplicator=>-5139, --- -0.313659667969 + j-0.949523925781
            im_multiplicator=>-15557
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(918),
            data_im_in=>first_stage_im_out(918),
            product_re_out=>mul_re_out(918),
            product_im_out=>mul_im_out(918)
        );

    UMUL_919 : complex_multiplier
    generic map(
            re_multiplicator=>-6455, --- -0.393981933594 + j-0.919067382812
            im_multiplicator=>-15058
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(919),
            data_im_in=>first_stage_im_out(919),
            product_re_out=>mul_re_out(919),
            product_im_out=>mul_im_out(919)
        );

    UMUL_920 : complex_multiplier
    generic map(
            re_multiplicator=>-7723, --- -0.471374511719 + j-0.881896972656
            im_multiplicator=>-14449
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(920),
            data_im_in=>first_stage_im_out(920),
            product_re_out=>mul_re_out(920),
            product_im_out=>mul_im_out(920)
        );

    UMUL_921 : complex_multiplier
    generic map(
            re_multiplicator=>-8934, --- -0.545288085938 + j-0.838195800781
            im_multiplicator=>-13733
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(921),
            data_im_in=>first_stage_im_out(921),
            product_re_out=>mul_re_out(921),
            product_im_out=>mul_im_out(921)
        );

    UMUL_922 : complex_multiplier
    generic map(
            re_multiplicator=>-10079, --- -0.615173339844 + j-0.788330078125
            im_multiplicator=>-12916
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(922),
            data_im_in=>first_stage_im_out(922),
            product_re_out=>mul_re_out(922),
            product_im_out=>mul_im_out(922)
        );

    UMUL_923 : complex_multiplier
    generic map(
            re_multiplicator=>-11150, --- -0.680541992188 + j-0.732604980469
            im_multiplicator=>-12003
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(923),
            data_im_in=>first_stage_im_out(923),
            product_re_out=>mul_re_out(923),
            product_im_out=>mul_im_out(923)
        );

    UMUL_924 : complex_multiplier
    generic map(
            re_multiplicator=>-12139, --- -0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(924),
            data_im_in=>first_stage_im_out(924),
            product_re_out=>mul_re_out(924),
            product_im_out=>mul_im_out(924)
        );

    UMUL_925 : complex_multiplier
    generic map(
            re_multiplicator=>-13038, --- -0.795776367188 + j-0.60546875
            im_multiplicator=>-9920
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(925),
            data_im_in=>first_stage_im_out(925),
            product_re_out=>mul_re_out(925),
            product_im_out=>mul_im_out(925)
        );

    UMUL_926 : complex_multiplier
    generic map(
            re_multiplicator=>-13842, --- -0.844848632812 + j-0.534973144531
            im_multiplicator=>-8765
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(926),
            data_im_in=>first_stage_im_out(926),
            product_re_out=>mul_re_out(926),
            product_im_out=>mul_im_out(926)
        );

    UMUL_927 : complex_multiplier
    generic map(
            re_multiplicator=>-14543, --- -0.887634277344 + j-0.460510253906
            im_multiplicator=>-7545
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(927),
            data_im_in=>first_stage_im_out(927),
            product_re_out=>mul_re_out(927),
            product_im_out=>mul_im_out(927)
        );

    UDELAY_928_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(928),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(928)
        );
    UDELAY_928_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(928),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(928)
        );
    USHIFTER_928_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(928),
            data_out=>mul_re_out(928)
        );
    USHIFTER_928_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(928),
            data_out=>mul_im_out(928)
        );

    UMUL_929 : complex_multiplier
    generic map(
            re_multiplicator=>16319, --- 0.996032714844 + j-0.0888061523438
            im_multiplicator=>-1455
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(929),
            data_im_in=>first_stage_im_out(929),
            product_re_out=>mul_re_out(929),
            product_im_out=>mul_im_out(929)
        );

    UMUL_930 : complex_multiplier
    generic map(
            re_multiplicator=>16125, --- 0.984191894531 + j-0.177001953125
            im_multiplicator=>-2900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(930),
            data_im_in=>first_stage_im_out(930),
            product_re_out=>mul_re_out(930),
            product_im_out=>mul_im_out(930)
        );

    UMUL_931 : complex_multiplier
    generic map(
            re_multiplicator=>15803, --- 0.964538574219 + j-0.263732910156
            im_multiplicator=>-4321
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(931),
            data_im_in=>first_stage_im_out(931),
            product_re_out=>mul_re_out(931),
            product_im_out=>mul_im_out(931)
        );

    UMUL_932 : complex_multiplier
    generic map(
            re_multiplicator=>15357, --- 0.937316894531 + j-0.348388671875
            im_multiplicator=>-5708
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(932),
            data_im_in=>first_stage_im_out(932),
            product_re_out=>mul_re_out(932),
            product_im_out=>mul_im_out(932)
        );

    UMUL_933 : complex_multiplier
    generic map(
            re_multiplicator=>14789, --- 0.902648925781 + j-0.430297851562
            im_multiplicator=>-7050
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(933),
            data_im_in=>first_stage_im_out(933),
            product_re_out=>mul_re_out(933),
            product_im_out=>mul_im_out(933)
        );

    UMUL_934 : complex_multiplier
    generic map(
            re_multiplicator=>14104, --- 0.86083984375 + j-0.5087890625
            im_multiplicator=>-8336
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(934),
            data_im_in=>first_stage_im_out(934),
            product_re_out=>mul_re_out(934),
            product_im_out=>mul_im_out(934)
        );

    UMUL_935 : complex_multiplier
    generic map(
            re_multiplicator=>13307, --- 0.812194824219 + j-0.583251953125
            im_multiplicator=>-9556
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(935),
            data_im_in=>first_stage_im_out(935),
            product_re_out=>mul_re_out(935),
            product_im_out=>mul_im_out(935)
        );

    UMUL_936 : complex_multiplier
    generic map(
            re_multiplicator=>12406, --- 0.757202148438 + j-0.653137207031
            im_multiplicator=>-10701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(936),
            data_im_in=>first_stage_im_out(936),
            product_re_out=>mul_re_out(936),
            product_im_out=>mul_im_out(936)
        );

    UMUL_937 : complex_multiplier
    generic map(
            re_multiplicator=>11406, --- 0.696166992188 + j-0.717834472656
            im_multiplicator=>-11761
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(937),
            data_im_in=>first_stage_im_out(937),
            product_re_out=>mul_re_out(937),
            product_im_out=>mul_im_out(937)
        );

    UMUL_938 : complex_multiplier
    generic map(
            re_multiplicator=>10315, --- 0.629577636719 + j-0.77685546875
            im_multiplicator=>-12728
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(938),
            data_im_in=>first_stage_im_out(938),
            product_re_out=>mul_re_out(938),
            product_im_out=>mul_im_out(938)
        );

    UMUL_939 : complex_multiplier
    generic map(
            re_multiplicator=>9144, --- 0.55810546875 + j-0.829711914062
            im_multiplicator=>-13594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(939),
            data_im_in=>first_stage_im_out(939),
            product_re_out=>mul_re_out(939),
            product_im_out=>mul_im_out(939)
        );

    UMUL_940 : complex_multiplier
    generic map(
            re_multiplicator=>7900, --- 0.482177734375 + j-0.876037597656
            im_multiplicator=>-14353
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(940),
            data_im_in=>first_stage_im_out(940),
            product_re_out=>mul_re_out(940),
            product_im_out=>mul_im_out(940)
        );

    UMUL_941 : complex_multiplier
    generic map(
            re_multiplicator=>6593, --- 0.402404785156 + j-0.915405273438
            im_multiplicator=>-14998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(941),
            data_im_in=>first_stage_im_out(941),
            product_re_out=>mul_re_out(941),
            product_im_out=>mul_im_out(941)
        );

    UMUL_942 : complex_multiplier
    generic map(
            re_multiplicator=>5234, --- 0.319458007812 + j-0.947570800781
            im_multiplicator=>-15525
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(942),
            data_im_in=>first_stage_im_out(942),
            product_re_out=>mul_re_out(942),
            product_im_out=>mul_im_out(942)
        );

    UMUL_943 : complex_multiplier
    generic map(
            re_multiplicator=>3834, --- 0.234008789062 + j-0.97216796875
            im_multiplicator=>-15928
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(943),
            data_im_in=>first_stage_im_out(943),
            product_re_out=>mul_re_out(943),
            product_im_out=>mul_im_out(943)
        );

    UMUL_944 : complex_multiplier
    generic map(
            re_multiplicator=>2404, --- 0.146728515625 + j-0.989135742188
            im_multiplicator=>-16206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(944),
            data_im_in=>first_stage_im_out(944),
            product_re_out=>mul_re_out(944),
            product_im_out=>mul_im_out(944)
        );

    UMUL_945 : complex_multiplier
    generic map(
            re_multiplicator=>954, --- 0.0582275390625 + j-0.998291015625
            im_multiplicator=>-16356
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(945),
            data_im_in=>first_stage_im_out(945),
            product_re_out=>mul_re_out(945),
            product_im_out=>mul_im_out(945)
        );

    UMUL_946 : complex_multiplier
    generic map(
            re_multiplicator=>-502, --- -0.0306396484375 + j-0.99951171875
            im_multiplicator=>-16376
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(946),
            data_im_in=>first_stage_im_out(946),
            product_re_out=>mul_re_out(946),
            product_im_out=>mul_im_out(946)
        );

    UMUL_947 : complex_multiplier
    generic map(
            re_multiplicator=>-1955, --- -0.119323730469 + j-0.992797851562
            im_multiplicator=>-16266
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(947),
            data_im_in=>first_stage_im_out(947),
            product_re_out=>mul_re_out(947),
            product_im_out=>mul_im_out(947)
        );

    UMUL_948 : complex_multiplier
    generic map(
            re_multiplicator=>-3393, --- -0.207092285156 + j-0.978271484375
            im_multiplicator=>-16028
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(948),
            data_im_in=>first_stage_im_out(948),
            product_re_out=>mul_re_out(948),
            product_im_out=>mul_im_out(948)
        );

    UMUL_949 : complex_multiplier
    generic map(
            re_multiplicator=>-4804, --- -0.293212890625 + j-0.955993652344
            im_multiplicator=>-15663
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(949),
            data_im_in=>first_stage_im_out(949),
            product_re_out=>mul_re_out(949),
            product_im_out=>mul_im_out(949)
        );

    UMUL_950 : complex_multiplier
    generic map(
            re_multiplicator=>-6176, --- -0.376953125 + j-0.926208496094
            im_multiplicator=>-15175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(950),
            data_im_in=>first_stage_im_out(950),
            product_re_out=>mul_re_out(950),
            product_im_out=>mul_im_out(950)
        );

    UMUL_951 : complex_multiplier
    generic map(
            re_multiplicator=>-7500, --- -0.457763671875 + j-0.889038085938
            im_multiplicator=>-14566
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(951),
            data_im_in=>first_stage_im_out(951),
            product_re_out=>mul_re_out(951),
            product_im_out=>mul_im_out(951)
        );

    UMUL_952 : complex_multiplier
    generic map(
            re_multiplicator=>-8765, --- -0.534973144531 + j-0.844848632812
            im_multiplicator=>-13842
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(952),
            data_im_in=>first_stage_im_out(952),
            product_re_out=>mul_re_out(952),
            product_im_out=>mul_im_out(952)
        );

    UMUL_953 : complex_multiplier
    generic map(
            re_multiplicator=>-9960, --- -0.60791015625 + j-0.7939453125
            im_multiplicator=>-13008
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(953),
            data_im_in=>first_stage_im_out(953),
            product_re_out=>mul_re_out(953),
            product_im_out=>mul_im_out(953)
        );

    UMUL_954 : complex_multiplier
    generic map(
            re_multiplicator=>-11077, --- -0.676086425781 + j-0.73681640625
            im_multiplicator=>-12072
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(954),
            data_im_in=>first_stage_im_out(954),
            product_re_out=>mul_re_out(954),
            product_im_out=>mul_im_out(954)
        );

    UMUL_955 : complex_multiplier
    generic map(
            re_multiplicator=>-12105, --- -0.738830566406 + j-0.673828125
            im_multiplicator=>-11040
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(955),
            data_im_in=>first_stage_im_out(955),
            product_re_out=>mul_re_out(955),
            product_im_out=>mul_im_out(955)
        );

    UMUL_956 : complex_multiplier
    generic map(
            re_multiplicator=>-13038, --- -0.795776367188 + j-0.60546875
            im_multiplicator=>-9920
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(956),
            data_im_in=>first_stage_im_out(956),
            product_re_out=>mul_re_out(956),
            product_im_out=>mul_im_out(956)
        );

    UMUL_957 : complex_multiplier
    generic map(
            re_multiplicator=>-13868, --- -0.846435546875 + j-0.532348632812
            im_multiplicator=>-8722
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(957),
            data_im_in=>first_stage_im_out(957),
            product_re_out=>mul_re_out(957),
            product_im_out=>mul_im_out(957)
        );

    UMUL_958 : complex_multiplier
    generic map(
            re_multiplicator=>-14589, --- -0.890441894531 + j-0.455078125
            im_multiplicator=>-7456
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(958),
            data_im_in=>first_stage_im_out(958),
            product_re_out=>mul_re_out(958),
            product_im_out=>mul_im_out(958)
        );

    UMUL_959 : complex_multiplier
    generic map(
            re_multiplicator=>-15193, --- -0.927307128906 + j-0.374145507812
            im_multiplicator=>-6130
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(959),
            data_im_in=>first_stage_im_out(959),
            product_re_out=>mul_re_out(959),
            product_im_out=>mul_im_out(959)
        );

    UDELAY_960_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(960),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(960)
        );
    UDELAY_960_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(960),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(960)
        );
    USHIFTER_960_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(960),
            data_out=>mul_re_out(960)
        );
    USHIFTER_960_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(960),
            data_out=>mul_im_out(960)
        );

    UMUL_961 : complex_multiplier
    generic map(
            re_multiplicator=>16314, --- 0.995727539062 + j-0.0918579101562
            im_multiplicator=>-1505
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(961),
            data_im_in=>first_stage_im_out(961),
            product_re_out=>mul_re_out(961),
            product_im_out=>mul_im_out(961)
        );

    UMUL_962 : complex_multiplier
    generic map(
            re_multiplicator=>16107, --- 0.983093261719 + j-0.182983398438
            im_multiplicator=>-2998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(962),
            data_im_in=>first_stage_im_out(962),
            product_re_out=>mul_re_out(962),
            product_im_out=>mul_im_out(962)
        );

    UMUL_963 : complex_multiplier
    generic map(
            re_multiplicator=>15763, --- 0.962097167969 + j-0.272583007812
            im_multiplicator=>-4466
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(963),
            data_im_in=>first_stage_im_out(963),
            product_re_out=>mul_re_out(963),
            product_im_out=>mul_im_out(963)
        );

    UMUL_964 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(964),
            data_im_in=>first_stage_im_out(964),
            product_re_out=>mul_re_out(964),
            product_im_out=>mul_im_out(964)
        );

    UMUL_965 : complex_multiplier
    generic map(
            re_multiplicator=>14679, --- 0.895935058594 + j-0.444091796875
            im_multiplicator=>-7276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(965),
            data_im_in=>first_stage_im_out(965),
            product_re_out=>mul_re_out(965),
            product_im_out=>mul_im_out(965)
        );

    UMUL_966 : complex_multiplier
    generic map(
            re_multiplicator=>13948, --- 0.851318359375 + j-0.524536132812
            im_multiplicator=>-8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(966),
            data_im_in=>first_stage_im_out(966),
            product_re_out=>mul_re_out(966),
            product_im_out=>mul_im_out(966)
        );

    UMUL_967 : complex_multiplier
    generic map(
            re_multiplicator=>13099, --- 0.799499511719 + j-0.6005859375
            im_multiplicator=>-9840
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(967),
            data_im_in=>first_stage_im_out(967),
            product_re_out=>mul_re_out(967),
            product_im_out=>mul_im_out(967)
        );

    UMUL_968 : complex_multiplier
    generic map(
            re_multiplicator=>12139, --- 0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(968),
            data_im_in=>first_stage_im_out(968),
            product_re_out=>mul_re_out(968),
            product_im_out=>mul_im_out(968)
        );

    UMUL_969 : complex_multiplier
    generic map(
            re_multiplicator=>11077, --- 0.676086425781 + j-0.73681640625
            im_multiplicator=>-12072
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(969),
            data_im_in=>first_stage_im_out(969),
            product_re_out=>mul_re_out(969),
            product_im_out=>mul_im_out(969)
        );

    UMUL_970 : complex_multiplier
    generic map(
            re_multiplicator=>9920, --- 0.60546875 + j-0.795776367188
            im_multiplicator=>-13038
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(970),
            data_im_in=>first_stage_im_out(970),
            product_re_out=>mul_re_out(970),
            product_im_out=>mul_im_out(970)
        );

    UMUL_971 : complex_multiplier
    generic map(
            re_multiplicator=>8680, --- 0.52978515625 + j-0.848083496094
            im_multiplicator=>-13895
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(971),
            data_im_in=>first_stage_im_out(971),
            product_re_out=>mul_re_out(971),
            product_im_out=>mul_im_out(971)
        );

    UMUL_972 : complex_multiplier
    generic map(
            re_multiplicator=>7366, --- 0.449584960938 + j-0.893188476562
            im_multiplicator=>-14634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(972),
            data_im_in=>first_stage_im_out(972),
            product_re_out=>mul_re_out(972),
            product_im_out=>mul_im_out(972)
        );

    UMUL_973 : complex_multiplier
    generic map(
            re_multiplicator=>5990, --- 0.365600585938 + j-0.930725097656
            im_multiplicator=>-15249
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(973),
            data_im_in=>first_stage_im_out(973),
            product_re_out=>mul_re_out(973),
            product_im_out=>mul_im_out(973)
        );

    UMUL_974 : complex_multiplier
    generic map(
            re_multiplicator=>4563, --- 0.278503417969 + j-0.960388183594
            im_multiplicator=>-15735
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(974),
            data_im_in=>first_stage_im_out(974),
            product_re_out=>mul_re_out(974),
            product_im_out=>mul_im_out(974)
        );

    UMUL_975 : complex_multiplier
    generic map(
            re_multiplicator=>3097, --- 0.189025878906 + j-0.98193359375
            im_multiplicator=>-16088
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(975),
            data_im_in=>first_stage_im_out(975),
            product_re_out=>mul_re_out(975),
            product_im_out=>mul_im_out(975)
        );

    UMUL_976 : complex_multiplier
    generic map(
            re_multiplicator=>1605, --- 0.0979614257812 + j-0.995178222656
            im_multiplicator=>-16305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(976),
            data_im_in=>first_stage_im_out(976),
            product_re_out=>mul_re_out(976),
            product_im_out=>mul_im_out(976)
        );

    UMUL_977 : complex_multiplier
    generic map(
            re_multiplicator=>100, --- 0.006103515625 + j-0.999938964844
            im_multiplicator=>-16383
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(977),
            data_im_in=>first_stage_im_out(977),
            product_re_out=>mul_re_out(977),
            product_im_out=>mul_im_out(977)
        );

    UMUL_978 : complex_multiplier
    generic map(
            re_multiplicator=>-1405, --- -0.0857543945312 + j-0.996276855469
            im_multiplicator=>-16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(978),
            data_im_in=>first_stage_im_out(978),
            product_re_out=>mul_re_out(978),
            product_im_out=>mul_im_out(978)
        );

    UMUL_979 : complex_multiplier
    generic map(
            re_multiplicator=>-2900, --- -0.177001953125 + j-0.984191894531
            im_multiplicator=>-16125
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(979),
            data_im_in=>first_stage_im_out(979),
            product_re_out=>mul_re_out(979),
            product_im_out=>mul_im_out(979)
        );

    UMUL_980 : complex_multiplier
    generic map(
            re_multiplicator=>-4369, --- -0.266662597656 + j-0.963745117188
            im_multiplicator=>-15790
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(980),
            data_im_in=>first_stage_im_out(980),
            product_re_out=>mul_re_out(980),
            product_im_out=>mul_im_out(980)
        );

    UMUL_981 : complex_multiplier
    generic map(
            re_multiplicator=>-5802, --- -0.354125976562 + j-0.935180664062
            im_multiplicator=>-15322
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(981),
            data_im_in=>first_stage_im_out(981),
            product_re_out=>mul_re_out(981),
            product_im_out=>mul_im_out(981)
        );

    UMUL_982 : complex_multiplier
    generic map(
            re_multiplicator=>-7186, --- -0.438598632812 + j-0.898620605469
            im_multiplicator=>-14723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(982),
            data_im_in=>first_stage_im_out(982),
            product_re_out=>mul_re_out(982),
            product_im_out=>mul_im_out(982)
        );

    UMUL_983 : complex_multiplier
    generic map(
            re_multiplicator=>-8509, --- -0.519348144531 + j-0.854553222656
            im_multiplicator=>-14001
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(983),
            data_im_in=>first_stage_im_out(983),
            product_re_out=>mul_re_out(983),
            product_im_out=>mul_im_out(983)
        );

    UMUL_984 : complex_multiplier
    generic map(
            re_multiplicator=>-9759, --- -0.595642089844 + j-0.803161621094
            im_multiplicator=>-13159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(984),
            data_im_in=>first_stage_im_out(984),
            product_re_out=>mul_re_out(984),
            product_im_out=>mul_im_out(984)
        );

    UMUL_985 : complex_multiplier
    generic map(
            re_multiplicator=>-10928, --- -0.6669921875 + j-0.745056152344
            im_multiplicator=>-12207
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(985),
            data_im_in=>first_stage_im_out(985),
            product_re_out=>mul_re_out(985),
            product_im_out=>mul_im_out(985)
        );

    UMUL_986 : complex_multiplier
    generic map(
            re_multiplicator=>-12003, --- -0.732604980469 + j-0.680541992188
            im_multiplicator=>-11150
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(986),
            data_im_in=>first_stage_im_out(986),
            product_re_out=>mul_re_out(986),
            product_im_out=>mul_im_out(986)
        );

    UMUL_987 : complex_multiplier
    generic map(
            re_multiplicator=>-12977, --- -0.792053222656 + j-0.6103515625
            im_multiplicator=>-10000
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(987),
            data_im_in=>first_stage_im_out(987),
            product_re_out=>mul_re_out(987),
            product_im_out=>mul_im_out(987)
        );

    UMUL_988 : complex_multiplier
    generic map(
            re_multiplicator=>-13842, --- -0.844848632812 + j-0.534973144531
            im_multiplicator=>-8765
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(988),
            data_im_in=>first_stage_im_out(988),
            product_re_out=>mul_re_out(988),
            product_im_out=>mul_im_out(988)
        );

    UMUL_989 : complex_multiplier
    generic map(
            re_multiplicator=>-14589, --- -0.890441894531 + j-0.455078125
            im_multiplicator=>-7456
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(989),
            data_im_in=>first_stage_im_out(989),
            product_re_out=>mul_re_out(989),
            product_im_out=>mul_im_out(989)
        );

    UMUL_990 : complex_multiplier
    generic map(
            re_multiplicator=>-15212, --- -0.928466796875 + j-0.371276855469
            im_multiplicator=>-6083
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(990),
            data_im_in=>first_stage_im_out(990),
            product_re_out=>mul_re_out(990),
            product_im_out=>mul_im_out(990)
        );

    UMUL_991 : complex_multiplier
    generic map(
            re_multiplicator=>-15707, --- -0.958679199219 + j-0.284362792969
            im_multiplicator=>-4659
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(991),
            data_im_in=>first_stage_im_out(991),
            product_re_out=>mul_re_out(991),
            product_im_out=>mul_im_out(991)
        );

    UDELAY_992_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(992),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(992)
        );
    UDELAY_992_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(992),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(992)
        );
    USHIFTER_992_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(992),
            data_out=>mul_re_out(992)
        );
    USHIFTER_992_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(992),
            data_out=>mul_im_out(992)
        );

    UMUL_993 : complex_multiplier
    generic map(
            re_multiplicator=>16309, --- 0.995422363281 + j-0.0949096679688
            im_multiplicator=>-1555
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(993),
            data_im_in=>first_stage_im_out(993),
            product_re_out=>mul_re_out(993),
            product_im_out=>mul_im_out(993)
        );

    UMUL_994 : complex_multiplier
    generic map(
            re_multiplicator=>16088, --- 0.98193359375 + j-0.189025878906
            im_multiplicator=>-3097
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(994),
            data_im_in=>first_stage_im_out(994),
            product_re_out=>mul_re_out(994),
            product_im_out=>mul_im_out(994)
        );

    UMUL_995 : complex_multiplier
    generic map(
            re_multiplicator=>15721, --- 0.959533691406 + j-0.281433105469
            im_multiplicator=>-4611
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(995),
            data_im_in=>first_stage_im_out(995),
            product_re_out=>mul_re_out(995),
            product_im_out=>mul_im_out(995)
        );

    UMUL_996 : complex_multiplier
    generic map(
            re_multiplicator=>15212, --- 0.928466796875 + j-0.371276855469
            im_multiplicator=>-6083
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(996),
            data_im_in=>first_stage_im_out(996),
            product_re_out=>mul_re_out(996),
            product_im_out=>mul_im_out(996)
        );

    UMUL_997 : complex_multiplier
    generic map(
            re_multiplicator=>14566, --- 0.889038085938 + j-0.457763671875
            im_multiplicator=>-7500
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(997),
            data_im_in=>first_stage_im_out(997),
            product_re_out=>mul_re_out(997),
            product_im_out=>mul_im_out(997)
        );

    UMUL_998 : complex_multiplier
    generic map(
            re_multiplicator=>13788, --- 0.841552734375 + j-0.540161132812
            im_multiplicator=>-8850
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(998),
            data_im_in=>first_stage_im_out(998),
            product_re_out=>mul_re_out(998),
            product_im_out=>mul_im_out(998)
        );

    UMUL_999 : complex_multiplier
    generic map(
            re_multiplicator=>12885, --- 0.786437988281 + j-0.617614746094
            im_multiplicator=>-10119
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(999),
            data_im_in=>first_stage_im_out(999),
            product_re_out=>mul_re_out(999),
            product_im_out=>mul_im_out(999)
        );

    UMUL_1000 : complex_multiplier
    generic map(
            re_multiplicator=>11866, --- 0.724243164062 + j-0.689514160156
            im_multiplicator=>-11297
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1000),
            data_im_in=>first_stage_im_out(1000),
            product_re_out=>mul_re_out(1000),
            product_im_out=>mul_im_out(1000)
        );

    UMUL_1001 : complex_multiplier
    generic map(
            re_multiplicator=>10739, --- 0.655456542969 + j-0.755187988281
            im_multiplicator=>-12373
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1001),
            data_im_in=>first_stage_im_out(1001),
            product_re_out=>mul_re_out(1001),
            product_im_out=>mul_im_out(1001)
        );

    UMUL_1002 : complex_multiplier
    generic map(
            re_multiplicator=>9516, --- 0.580810546875 + j-0.814025878906
            im_multiplicator=>-13337
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1002),
            data_im_in=>first_stage_im_out(1002),
            product_re_out=>mul_re_out(1002),
            product_im_out=>mul_im_out(1002)
        );

    UMUL_1003 : complex_multiplier
    generic map(
            re_multiplicator=>8206, --- 0.500854492188 + j-0.865478515625
            im_multiplicator=>-14180
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1003),
            data_im_in=>first_stage_im_out(1003),
            product_re_out=>mul_re_out(1003),
            product_im_out=>mul_im_out(1003)
        );

    UMUL_1004 : complex_multiplier
    generic map(
            re_multiplicator=>6822, --- 0.416381835938 + j-0.909118652344
            im_multiplicator=>-14895
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1004),
            data_im_in=>first_stage_im_out(1004),
            product_re_out=>mul_re_out(1004),
            product_im_out=>mul_im_out(1004)
        );

    UMUL_1005 : complex_multiplier
    generic map(
            re_multiplicator=>5377, --- 0.328186035156 + j-0.944580078125
            im_multiplicator=>-15476
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1005),
            data_im_in=>first_stage_im_out(1005),
            product_re_out=>mul_re_out(1005),
            product_im_out=>mul_im_out(1005)
        );

    UMUL_1006 : complex_multiplier
    generic map(
            re_multiplicator=>3883, --- 0.236999511719 + j-0.971496582031
            im_multiplicator=>-15917
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1006),
            data_im_in=>first_stage_im_out(1006),
            product_re_out=>mul_re_out(1006),
            product_im_out=>mul_im_out(1006)
        );

    UMUL_1007 : complex_multiplier
    generic map(
            re_multiplicator=>2354, --- 0.143676757812 + j-0.989562988281
            im_multiplicator=>-16213
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1007),
            data_im_in=>first_stage_im_out(1007),
            product_re_out=>mul_re_out(1007),
            product_im_out=>mul_im_out(1007)
        );

    UMUL_1008 : complex_multiplier
    generic map(
            re_multiplicator=>803, --- 0.0490112304688 + j-0.998779296875
            im_multiplicator=>-16364
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1008),
            data_im_in=>first_stage_im_out(1008),
            product_re_out=>mul_re_out(1008),
            product_im_out=>mul_im_out(1008)
        );

    UMUL_1009 : complex_multiplier
    generic map(
            re_multiplicator=>-753, --- -0.0459594726562 + j-0.998901367188
            im_multiplicator=>-16366
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1009),
            data_im_in=>first_stage_im_out(1009),
            product_re_out=>mul_re_out(1009),
            product_im_out=>mul_im_out(1009)
        );

    UMUL_1010 : complex_multiplier
    generic map(
            re_multiplicator=>-2304, --- -0.140625 + j-0.990051269531
            im_multiplicator=>-16221
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1010),
            data_im_in=>first_stage_im_out(1010),
            product_re_out=>mul_re_out(1010),
            product_im_out=>mul_im_out(1010)
        );

    UMUL_1011 : complex_multiplier
    generic map(
            re_multiplicator=>-3834, --- -0.234008789062 + j-0.97216796875
            im_multiplicator=>-15928
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1011),
            data_im_in=>first_stage_im_out(1011),
            product_re_out=>mul_re_out(1011),
            product_im_out=>mul_im_out(1011)
        );

    UMUL_1012 : complex_multiplier
    generic map(
            re_multiplicator=>-5329, --- -0.325256347656 + j-0.945556640625
            im_multiplicator=>-15492
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1012),
            data_im_in=>first_stage_im_out(1012),
            product_re_out=>mul_re_out(1012),
            product_im_out=>mul_im_out(1012)
        );

    UMUL_1013 : complex_multiplier
    generic map(
            re_multiplicator=>-6777, --- -0.413635253906 + j-0.910400390625
            im_multiplicator=>-14916
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1013),
            data_im_in=>first_stage_im_out(1013),
            product_re_out=>mul_re_out(1013),
            product_im_out=>mul_im_out(1013)
        );

    UMUL_1014 : complex_multiplier
    generic map(
            re_multiplicator=>-8162, --- -0.498168945312 + j-0.867004394531
            im_multiplicator=>-14205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1014),
            data_im_in=>first_stage_im_out(1014),
            product_re_out=>mul_re_out(1014),
            product_im_out=>mul_im_out(1014)
        );

    UMUL_1015 : complex_multiplier
    generic map(
            re_multiplicator=>-9475, --- -0.578308105469 + j-0.815795898438
            im_multiplicator=>-13366
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1015),
            data_im_in=>first_stage_im_out(1015),
            product_re_out=>mul_re_out(1015),
            product_im_out=>mul_im_out(1015)
        );

    UMUL_1016 : complex_multiplier
    generic map(
            re_multiplicator=>-10701, --- -0.653137207031 + j-0.757202148438
            im_multiplicator=>-12406
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1016),
            data_im_in=>first_stage_im_out(1016),
            product_re_out=>mul_re_out(1016),
            product_im_out=>mul_im_out(1016)
        );

    UMUL_1017 : complex_multiplier
    generic map(
            re_multiplicator=>-11831, --- -0.722106933594 + j-0.691711425781
            im_multiplicator=>-11333
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1017),
            data_im_in=>first_stage_im_out(1017),
            product_re_out=>mul_re_out(1017),
            product_im_out=>mul_im_out(1017)
        );

    UMUL_1018 : complex_multiplier
    generic map(
            re_multiplicator=>-12854, --- -0.784545898438 + j-0.620056152344
            im_multiplicator=>-10159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1018),
            data_im_in=>first_stage_im_out(1018),
            product_re_out=>mul_re_out(1018),
            product_im_out=>mul_im_out(1018)
        );

    UMUL_1019 : complex_multiplier
    generic map(
            re_multiplicator=>-13760, --- -0.83984375 + j-0.542724609375
            im_multiplicator=>-8892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1019),
            data_im_in=>first_stage_im_out(1019),
            product_re_out=>mul_re_out(1019),
            product_im_out=>mul_im_out(1019)
        );

    UMUL_1020 : complex_multiplier
    generic map(
            re_multiplicator=>-14543, --- -0.887634277344 + j-0.460510253906
            im_multiplicator=>-7545
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1020),
            data_im_in=>first_stage_im_out(1020),
            product_re_out=>mul_re_out(1020),
            product_im_out=>mul_im_out(1020)
        );

    UMUL_1021 : complex_multiplier
    generic map(
            re_multiplicator=>-15193, --- -0.927307128906 + j-0.374145507812
            im_multiplicator=>-6130
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1021),
            data_im_in=>first_stage_im_out(1021),
            product_re_out=>mul_re_out(1021),
            product_im_out=>mul_im_out(1021)
        );

    UMUL_1022 : complex_multiplier
    generic map(
            re_multiplicator=>-15707, --- -0.958679199219 + j-0.284362792969
            im_multiplicator=>-4659
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1022),
            data_im_in=>first_stage_im_out(1022),
            product_re_out=>mul_re_out(1022),
            product_im_out=>mul_im_out(1022)
        );

    UMUL_1023 : complex_multiplier
    generic map(
            re_multiplicator=>-16078, --- -0.981323242188 + j-0.192077636719
            im_multiplicator=>-3147
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1023),
            data_im_in=>first_stage_im_out(1023),
            product_re_out=>mul_re_out(1023),
            product_im_out=>mul_im_out(1023)
        );

    UDELAY_1024_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1024),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1024)
        );
    UDELAY_1024_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1024),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1024)
        );
    USHIFTER_1024_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1024),
            data_out=>mul_re_out(1024)
        );
    USHIFTER_1024_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1024),
            data_out=>mul_im_out(1024)
        );

    UMUL_1025 : complex_multiplier
    generic map(
            re_multiplicator=>16305, --- 0.995178222656 + j-0.0979614257812
            im_multiplicator=>-1605
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1025),
            data_im_in=>first_stage_im_out(1025),
            product_re_out=>mul_re_out(1025),
            product_im_out=>mul_im_out(1025)
        );

    UMUL_1026 : complex_multiplier
    generic map(
            re_multiplicator=>16069, --- 0.980773925781 + j-0.195068359375
            im_multiplicator=>-3196
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1026),
            data_im_in=>first_stage_im_out(1026),
            product_re_out=>mul_re_out(1026),
            product_im_out=>mul_im_out(1026)
        );

    UMUL_1027 : complex_multiplier
    generic map(
            re_multiplicator=>15678, --- 0.956909179688 + j-0.290283203125
            im_multiplicator=>-4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1027),
            data_im_in=>first_stage_im_out(1027),
            product_re_out=>mul_re_out(1027),
            product_im_out=>mul_im_out(1027)
        );

    UMUL_1028 : complex_multiplier
    generic map(
            re_multiplicator=>15136, --- 0.923828125 + j-0.382629394531
            im_multiplicator=>-6269
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1028),
            data_im_in=>first_stage_im_out(1028),
            product_re_out=>mul_re_out(1028),
            product_im_out=>mul_im_out(1028)
        );

    UMUL_1029 : complex_multiplier
    generic map(
            re_multiplicator=>14449, --- 0.881896972656 + j-0.471374511719
            im_multiplicator=>-7723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1029),
            data_im_in=>first_stage_im_out(1029),
            product_re_out=>mul_re_out(1029),
            product_im_out=>mul_im_out(1029)
        );

    UMUL_1030 : complex_multiplier
    generic map(
            re_multiplicator=>13622, --- 0.831420898438 + j-0.555541992188
            im_multiplicator=>-9102
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1030),
            data_im_in=>first_stage_im_out(1030),
            product_re_out=>mul_re_out(1030),
            product_im_out=>mul_im_out(1030)
        );

    UMUL_1031 : complex_multiplier
    generic map(
            re_multiplicator=>12665, --- 0.773010253906 + j-0.634338378906
            im_multiplicator=>-10393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1031),
            data_im_in=>first_stage_im_out(1031),
            product_re_out=>mul_re_out(1031),
            product_im_out=>mul_im_out(1031)
        );

    UMUL_1032 : complex_multiplier
    generic map(
            re_multiplicator=>11585, --- 0.707092285156 + j-0.707092285156
            im_multiplicator=>-11585
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1032),
            data_im_in=>first_stage_im_out(1032),
            product_re_out=>mul_re_out(1032),
            product_im_out=>mul_im_out(1032)
        );

    UMUL_1033 : complex_multiplier
    generic map(
            re_multiplicator=>10393, --- 0.634338378906 + j-0.773010253906
            im_multiplicator=>-12665
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1033),
            data_im_in=>first_stage_im_out(1033),
            product_re_out=>mul_re_out(1033),
            product_im_out=>mul_im_out(1033)
        );

    UMUL_1034 : complex_multiplier
    generic map(
            re_multiplicator=>9102, --- 0.555541992188 + j-0.831420898438
            im_multiplicator=>-13622
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1034),
            data_im_in=>first_stage_im_out(1034),
            product_re_out=>mul_re_out(1034),
            product_im_out=>mul_im_out(1034)
        );

    UMUL_1035 : complex_multiplier
    generic map(
            re_multiplicator=>7723, --- 0.471374511719 + j-0.881896972656
            im_multiplicator=>-14449
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1035),
            data_im_in=>first_stage_im_out(1035),
            product_re_out=>mul_re_out(1035),
            product_im_out=>mul_im_out(1035)
        );

    UMUL_1036 : complex_multiplier
    generic map(
            re_multiplicator=>6269, --- 0.382629394531 + j-0.923828125
            im_multiplicator=>-15136
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1036),
            data_im_in=>first_stage_im_out(1036),
            product_re_out=>mul_re_out(1036),
            product_im_out=>mul_im_out(1036)
        );

    UMUL_1037 : complex_multiplier
    generic map(
            re_multiplicator=>4756, --- 0.290283203125 + j-0.956909179688
            im_multiplicator=>-15678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1037),
            data_im_in=>first_stage_im_out(1037),
            product_re_out=>mul_re_out(1037),
            product_im_out=>mul_im_out(1037)
        );

    UMUL_1038 : complex_multiplier
    generic map(
            re_multiplicator=>3196, --- 0.195068359375 + j-0.980773925781
            im_multiplicator=>-16069
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1038),
            data_im_in=>first_stage_im_out(1038),
            product_re_out=>mul_re_out(1038),
            product_im_out=>mul_im_out(1038)
        );

    UMUL_1039 : complex_multiplier
    generic map(
            re_multiplicator=>1605, --- 0.0979614257812 + j-0.995178222656
            im_multiplicator=>-16305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1039),
            data_im_in=>first_stage_im_out(1039),
            product_re_out=>mul_re_out(1039),
            product_im_out=>mul_im_out(1039)
        );

    UMUL_1040 : complex_multiplier
    generic map(
            re_multiplicator=>0, --- 0.0 + j-1.0
            im_multiplicator=>-16384
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1040),
            data_im_in=>first_stage_im_out(1040),
            product_re_out=>mul_re_out(1040),
            product_im_out=>mul_im_out(1040)
        );

    UMUL_1041 : complex_multiplier
    generic map(
            re_multiplicator=>-1605, --- -0.0979614257812 + j-0.995178222656
            im_multiplicator=>-16305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1041),
            data_im_in=>first_stage_im_out(1041),
            product_re_out=>mul_re_out(1041),
            product_im_out=>mul_im_out(1041)
        );

    UMUL_1042 : complex_multiplier
    generic map(
            re_multiplicator=>-3196, --- -0.195068359375 + j-0.980773925781
            im_multiplicator=>-16069
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1042),
            data_im_in=>first_stage_im_out(1042),
            product_re_out=>mul_re_out(1042),
            product_im_out=>mul_im_out(1042)
        );

    UMUL_1043 : complex_multiplier
    generic map(
            re_multiplicator=>-4756, --- -0.290283203125 + j-0.956909179688
            im_multiplicator=>-15678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1043),
            data_im_in=>first_stage_im_out(1043),
            product_re_out=>mul_re_out(1043),
            product_im_out=>mul_im_out(1043)
        );

    UMUL_1044 : complex_multiplier
    generic map(
            re_multiplicator=>-6269, --- -0.382629394531 + j-0.923828125
            im_multiplicator=>-15136
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1044),
            data_im_in=>first_stage_im_out(1044),
            product_re_out=>mul_re_out(1044),
            product_im_out=>mul_im_out(1044)
        );

    UMUL_1045 : complex_multiplier
    generic map(
            re_multiplicator=>-7723, --- -0.471374511719 + j-0.881896972656
            im_multiplicator=>-14449
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1045),
            data_im_in=>first_stage_im_out(1045),
            product_re_out=>mul_re_out(1045),
            product_im_out=>mul_im_out(1045)
        );

    UMUL_1046 : complex_multiplier
    generic map(
            re_multiplicator=>-9102, --- -0.555541992188 + j-0.831420898438
            im_multiplicator=>-13622
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1046),
            data_im_in=>first_stage_im_out(1046),
            product_re_out=>mul_re_out(1046),
            product_im_out=>mul_im_out(1046)
        );

    UMUL_1047 : complex_multiplier
    generic map(
            re_multiplicator=>-10393, --- -0.634338378906 + j-0.773010253906
            im_multiplicator=>-12665
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1047),
            data_im_in=>first_stage_im_out(1047),
            product_re_out=>mul_re_out(1047),
            product_im_out=>mul_im_out(1047)
        );

    UMUL_1048 : complex_multiplier
    generic map(
            re_multiplicator=>-11585, --- -0.707092285156 + j-0.707092285156
            im_multiplicator=>-11585
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1048),
            data_im_in=>first_stage_im_out(1048),
            product_re_out=>mul_re_out(1048),
            product_im_out=>mul_im_out(1048)
        );

    UMUL_1049 : complex_multiplier
    generic map(
            re_multiplicator=>-12665, --- -0.773010253906 + j-0.634338378906
            im_multiplicator=>-10393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1049),
            data_im_in=>first_stage_im_out(1049),
            product_re_out=>mul_re_out(1049),
            product_im_out=>mul_im_out(1049)
        );

    UMUL_1050 : complex_multiplier
    generic map(
            re_multiplicator=>-13622, --- -0.831420898438 + j-0.555541992188
            im_multiplicator=>-9102
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1050),
            data_im_in=>first_stage_im_out(1050),
            product_re_out=>mul_re_out(1050),
            product_im_out=>mul_im_out(1050)
        );

    UMUL_1051 : complex_multiplier
    generic map(
            re_multiplicator=>-14449, --- -0.881896972656 + j-0.471374511719
            im_multiplicator=>-7723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1051),
            data_im_in=>first_stage_im_out(1051),
            product_re_out=>mul_re_out(1051),
            product_im_out=>mul_im_out(1051)
        );

    UMUL_1052 : complex_multiplier
    generic map(
            re_multiplicator=>-15136, --- -0.923828125 + j-0.382629394531
            im_multiplicator=>-6269
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1052),
            data_im_in=>first_stage_im_out(1052),
            product_re_out=>mul_re_out(1052),
            product_im_out=>mul_im_out(1052)
        );

    UMUL_1053 : complex_multiplier
    generic map(
            re_multiplicator=>-15678, --- -0.956909179688 + j-0.290283203125
            im_multiplicator=>-4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1053),
            data_im_in=>first_stage_im_out(1053),
            product_re_out=>mul_re_out(1053),
            product_im_out=>mul_im_out(1053)
        );

    UMUL_1054 : complex_multiplier
    generic map(
            re_multiplicator=>-16069, --- -0.980773925781 + j-0.195068359375
            im_multiplicator=>-3196
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1054),
            data_im_in=>first_stage_im_out(1054),
            product_re_out=>mul_re_out(1054),
            product_im_out=>mul_im_out(1054)
        );

    UMUL_1055 : complex_multiplier
    generic map(
            re_multiplicator=>-16305, --- -0.995178222656 + j-0.0979614257812
            im_multiplicator=>-1605
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1055),
            data_im_in=>first_stage_im_out(1055),
            product_re_out=>mul_re_out(1055),
            product_im_out=>mul_im_out(1055)
        );

    UDELAY_1056_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1056),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1056)
        );
    UDELAY_1056_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1056),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1056)
        );
    USHIFTER_1056_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1056),
            data_out=>mul_re_out(1056)
        );
    USHIFTER_1056_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1056),
            data_out=>mul_im_out(1056)
        );

    UMUL_1057 : complex_multiplier
    generic map(
            re_multiplicator=>16300, --- 0.994873046875 + j-0.101013183594
            im_multiplicator=>-1655
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1057),
            data_im_in=>first_stage_im_out(1057),
            product_re_out=>mul_re_out(1057),
            product_im_out=>mul_im_out(1057)
        );

    UMUL_1058 : complex_multiplier
    generic map(
            re_multiplicator=>16049, --- 0.979553222656 + j-0.201049804688
            im_multiplicator=>-3294
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1058),
            data_im_in=>first_stage_im_out(1058),
            product_re_out=>mul_re_out(1058),
            product_im_out=>mul_im_out(1058)
        );

    UMUL_1059 : complex_multiplier
    generic map(
            re_multiplicator=>15634, --- 0.954223632812 + j-0.299072265625
            im_multiplicator=>-4900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1059),
            data_im_in=>first_stage_im_out(1059),
            product_re_out=>mul_re_out(1059),
            product_im_out=>mul_im_out(1059)
        );

    UMUL_1060 : complex_multiplier
    generic map(
            re_multiplicator=>15058, --- 0.919067382812 + j-0.393981933594
            im_multiplicator=>-6455
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1060),
            data_im_in=>first_stage_im_out(1060),
            product_re_out=>mul_re_out(1060),
            product_im_out=>mul_im_out(1060)
        );

    UMUL_1061 : complex_multiplier
    generic map(
            re_multiplicator=>14329, --- 0.874572753906 + j-0.48486328125
            im_multiplicator=>-7944
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1061),
            data_im_in=>first_stage_im_out(1061),
            product_re_out=>mul_re_out(1061),
            product_im_out=>mul_im_out(1061)
        );

    UMUL_1062 : complex_multiplier
    generic map(
            re_multiplicator=>13452, --- 0.821044921875 + j-0.570739746094
            im_multiplicator=>-9351
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1062),
            data_im_in=>first_stage_im_out(1062),
            product_re_out=>mul_re_out(1062),
            product_im_out=>mul_im_out(1062)
        );

    UMUL_1063 : complex_multiplier
    generic map(
            re_multiplicator=>12438, --- 0.759155273438 + j-0.650817871094
            im_multiplicator=>-10663
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1063),
            data_im_in=>first_stage_im_out(1063),
            product_re_out=>mul_re_out(1063),
            product_im_out=>mul_im_out(1063)
        );

    UMUL_1064 : complex_multiplier
    generic map(
            re_multiplicator=>11297, --- 0.689514160156 + j-0.724243164062
            im_multiplicator=>-11866
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1064),
            data_im_in=>first_stage_im_out(1064),
            product_re_out=>mul_re_out(1064),
            product_im_out=>mul_im_out(1064)
        );

    UMUL_1065 : complex_multiplier
    generic map(
            re_multiplicator=>10040, --- 0.61279296875 + j-0.790222167969
            im_multiplicator=>-12947
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1065),
            data_im_in=>first_stage_im_out(1065),
            product_re_out=>mul_re_out(1065),
            product_im_out=>mul_im_out(1065)
        );

    UMUL_1066 : complex_multiplier
    generic map(
            re_multiplicator=>8680, --- 0.52978515625 + j-0.848083496094
            im_multiplicator=>-13895
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1066),
            data_im_in=>first_stage_im_out(1066),
            product_re_out=>mul_re_out(1066),
            product_im_out=>mul_im_out(1066)
        );

    UMUL_1067 : complex_multiplier
    generic map(
            re_multiplicator=>7231, --- 0.441345214844 + j-0.897277832031
            im_multiplicator=>-14701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1067),
            data_im_in=>first_stage_im_out(1067),
            product_re_out=>mul_re_out(1067),
            product_im_out=>mul_im_out(1067)
        );

    UMUL_1068 : complex_multiplier
    generic map(
            re_multiplicator=>5708, --- 0.348388671875 + j-0.937316894531
            im_multiplicator=>-15357
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1068),
            data_im_in=>first_stage_im_out(1068),
            product_re_out=>mul_re_out(1068),
            product_im_out=>mul_im_out(1068)
        );

    UMUL_1069 : complex_multiplier
    generic map(
            re_multiplicator=>4127, --- 0.251892089844 + j-0.967712402344
            im_multiplicator=>-15855
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1069),
            data_im_in=>first_stage_im_out(1069),
            product_re_out=>mul_re_out(1069),
            product_im_out=>mul_im_out(1069)
        );

    UMUL_1070 : complex_multiplier
    generic map(
            re_multiplicator=>2503, --- 0.152770996094 + j-0.988220214844
            im_multiplicator=>-16191
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1070),
            data_im_in=>first_stage_im_out(1070),
            product_re_out=>mul_re_out(1070),
            product_im_out=>mul_im_out(1070)
        );

    UMUL_1071 : complex_multiplier
    generic map(
            re_multiplicator=>854, --- 0.0521240234375 + j-0.998596191406
            im_multiplicator=>-16361
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1071),
            data_im_in=>first_stage_im_out(1071),
            product_re_out=>mul_re_out(1071),
            product_im_out=>mul_im_out(1071)
        );

    UMUL_1072 : complex_multiplier
    generic map(
            re_multiplicator=>-803, --- -0.0490112304688 + j-0.998779296875
            im_multiplicator=>-16364
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1072),
            data_im_in=>first_stage_im_out(1072),
            product_re_out=>mul_re_out(1072),
            product_im_out=>mul_im_out(1072)
        );

    UMUL_1073 : complex_multiplier
    generic map(
            re_multiplicator=>-2453, --- -0.149719238281 + j-0.988708496094
            im_multiplicator=>-16199
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1073),
            data_im_in=>first_stage_im_out(1073),
            product_re_out=>mul_re_out(1073),
            product_im_out=>mul_im_out(1073)
        );

    UMUL_1074 : complex_multiplier
    generic map(
            re_multiplicator=>-4078, --- -0.248901367188 + j-0.968505859375
            im_multiplicator=>-15868
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1074),
            data_im_in=>first_stage_im_out(1074),
            product_re_out=>mul_re_out(1074),
            product_im_out=>mul_im_out(1074)
        );

    UMUL_1075 : complex_multiplier
    generic map(
            re_multiplicator=>-5661, --- -0.345520019531 + j-0.938354492188
            im_multiplicator=>-15374
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1075),
            data_im_in=>first_stage_im_out(1075),
            product_re_out=>mul_re_out(1075),
            product_im_out=>mul_im_out(1075)
        );

    UMUL_1076 : complex_multiplier
    generic map(
            re_multiplicator=>-7186, --- -0.438598632812 + j-0.898620605469
            im_multiplicator=>-14723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1076),
            data_im_in=>first_stage_im_out(1076),
            product_re_out=>mul_re_out(1076),
            product_im_out=>mul_im_out(1076)
        );

    UMUL_1077 : complex_multiplier
    generic map(
            re_multiplicator=>-8637, --- -0.527160644531 + j-0.849731445312
            im_multiplicator=>-13922
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1077),
            data_im_in=>first_stage_im_out(1077),
            product_re_out=>mul_re_out(1077),
            product_im_out=>mul_im_out(1077)
        );

    UMUL_1078 : complex_multiplier
    generic map(
            re_multiplicator=>-10000, --- -0.6103515625 + j-0.792053222656
            im_multiplicator=>-12977
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1078),
            data_im_in=>first_stage_im_out(1078),
            product_re_out=>mul_re_out(1078),
            product_im_out=>mul_im_out(1078)
        );

    UMUL_1079 : complex_multiplier
    generic map(
            re_multiplicator=>-11260, --- -0.687255859375 + j-0.726318359375
            im_multiplicator=>-11900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1079),
            data_im_in=>first_stage_im_out(1079),
            product_re_out=>mul_re_out(1079),
            product_im_out=>mul_im_out(1079)
        );

    UMUL_1080 : complex_multiplier
    generic map(
            re_multiplicator=>-12406, --- -0.757202148438 + j-0.653137207031
            im_multiplicator=>-10701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1080),
            data_im_in=>first_stage_im_out(1080),
            product_re_out=>mul_re_out(1080),
            product_im_out=>mul_im_out(1080)
        );

    UMUL_1081 : complex_multiplier
    generic map(
            re_multiplicator=>-13424, --- -0.8193359375 + j-0.5732421875
            im_multiplicator=>-9392
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1081),
            data_im_in=>first_stage_im_out(1081),
            product_re_out=>mul_re_out(1081),
            product_im_out=>mul_im_out(1081)
        );

    UMUL_1082 : complex_multiplier
    generic map(
            re_multiplicator=>-14304, --- -0.873046875 + j-0.487548828125
            im_multiplicator=>-7988
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1082),
            data_im_in=>first_stage_im_out(1082),
            product_re_out=>mul_re_out(1082),
            product_im_out=>mul_im_out(1082)
        );

    UMUL_1083 : complex_multiplier
    generic map(
            re_multiplicator=>-15038, --- -0.917846679688 + j-0.396789550781
            im_multiplicator=>-6501
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1083),
            data_im_in=>first_stage_im_out(1083),
            product_re_out=>mul_re_out(1083),
            product_im_out=>mul_im_out(1083)
        );

    UMUL_1084 : complex_multiplier
    generic map(
            re_multiplicator=>-15618, --- -0.953247070312 + j-0.302001953125
            im_multiplicator=>-4948
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1084),
            data_im_in=>first_stage_im_out(1084),
            product_re_out=>mul_re_out(1084),
            product_im_out=>mul_im_out(1084)
        );

    UMUL_1085 : complex_multiplier
    generic map(
            re_multiplicator=>-16039, --- -0.978942871094 + j-0.2041015625
            im_multiplicator=>-3344
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1085),
            data_im_in=>first_stage_im_out(1085),
            product_re_out=>mul_re_out(1085),
            product_im_out=>mul_im_out(1085)
        );

    UMUL_1086 : complex_multiplier
    generic map(
            re_multiplicator=>-16294, --- -0.994506835938 + j-0.104064941406
            im_multiplicator=>-1705
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1086),
            data_im_in=>first_stage_im_out(1086),
            product_re_out=>mul_re_out(1086),
            product_im_out=>mul_im_out(1086)
        );

    UMUL_1087 : complex_multiplier
    generic map(
            re_multiplicator=>-16383, --- -0.999938964844 + j-0.0030517578125
            im_multiplicator=>-50
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1087),
            data_im_in=>first_stage_im_out(1087),
            product_re_out=>mul_re_out(1087),
            product_im_out=>mul_im_out(1087)
        );

    UDELAY_1088_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1088),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1088)
        );
    UDELAY_1088_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1088),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1088)
        );
    USHIFTER_1088_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1088),
            data_out=>mul_re_out(1088)
        );
    USHIFTER_1088_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1088),
            data_out=>mul_im_out(1088)
        );

    UMUL_1089 : complex_multiplier
    generic map(
            re_multiplicator=>16294, --- 0.994506835938 + j-0.104064941406
            im_multiplicator=>-1705
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1089),
            data_im_in=>first_stage_im_out(1089),
            product_re_out=>mul_re_out(1089),
            product_im_out=>mul_im_out(1089)
        );

    UMUL_1090 : complex_multiplier
    generic map(
            re_multiplicator=>16028, --- 0.978271484375 + j-0.207092285156
            im_multiplicator=>-3393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1090),
            data_im_in=>first_stage_im_out(1090),
            product_re_out=>mul_re_out(1090),
            product_im_out=>mul_im_out(1090)
        );

    UMUL_1091 : complex_multiplier
    generic map(
            re_multiplicator=>15588, --- 0.951416015625 + j-0.307800292969
            im_multiplicator=>-5043
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1091),
            data_im_in=>first_stage_im_out(1091),
            product_re_out=>mul_re_out(1091),
            product_im_out=>mul_im_out(1091)
        );

    UMUL_1092 : complex_multiplier
    generic map(
            re_multiplicator=>14978, --- 0.914184570312 + j-0.405212402344
            im_multiplicator=>-6639
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1092),
            data_im_in=>first_stage_im_out(1092),
            product_re_out=>mul_re_out(1092),
            product_im_out=>mul_im_out(1092)
        );

    UMUL_1093 : complex_multiplier
    generic map(
            re_multiplicator=>14205, --- 0.867004394531 + j-0.498168945312
            im_multiplicator=>-8162
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1093),
            data_im_in=>first_stage_im_out(1093),
            product_re_out=>mul_re_out(1093),
            product_im_out=>mul_im_out(1093)
        );

    UMUL_1094 : complex_multiplier
    generic map(
            re_multiplicator=>13278, --- 0.810424804688 + j-0.585754394531
            im_multiplicator=>-9597
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1094),
            data_im_in=>first_stage_im_out(1094),
            product_re_out=>mul_re_out(1094),
            product_im_out=>mul_im_out(1094)
        );

    UMUL_1095 : complex_multiplier
    generic map(
            re_multiplicator=>12207, --- 0.745056152344 + j-0.6669921875
            im_multiplicator=>-10928
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1095),
            data_im_in=>first_stage_im_out(1095),
            product_re_out=>mul_re_out(1095),
            product_im_out=>mul_im_out(1095)
        );

    UMUL_1096 : complex_multiplier
    generic map(
            re_multiplicator=>11002, --- 0.671508789062 + j-0.740905761719
            im_multiplicator=>-12139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1096),
            data_im_in=>first_stage_im_out(1096),
            product_re_out=>mul_re_out(1096),
            product_im_out=>mul_im_out(1096)
        );

    UMUL_1097 : complex_multiplier
    generic map(
            re_multiplicator=>9679, --- 0.590759277344 + j-0.806823730469
            im_multiplicator=>-13219
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1097),
            data_im_in=>first_stage_im_out(1097),
            product_re_out=>mul_re_out(1097),
            product_im_out=>mul_im_out(1097)
        );

    UMUL_1098 : complex_multiplier
    generic map(
            re_multiplicator=>8249, --- 0.503479003906 + j-0.863952636719
            im_multiplicator=>-14155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1098),
            data_im_in=>first_stage_im_out(1098),
            product_re_out=>mul_re_out(1098),
            product_im_out=>mul_im_out(1098)
        );

    UMUL_1099 : complex_multiplier
    generic map(
            re_multiplicator=>6731, --- 0.410827636719 + j-0.911682128906
            im_multiplicator=>-14937
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1099),
            data_im_in=>first_stage_im_out(1099),
            product_re_out=>mul_re_out(1099),
            product_im_out=>mul_im_out(1099)
        );

    UMUL_1100 : complex_multiplier
    generic map(
            re_multiplicator=>5139, --- 0.313659667969 + j-0.949523925781
            im_multiplicator=>-15557
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1100),
            data_im_in=>first_stage_im_out(1100),
            product_re_out=>mul_re_out(1100),
            product_im_out=>mul_im_out(1100)
        );

    UMUL_1101 : complex_multiplier
    generic map(
            re_multiplicator=>3491, --- 0.213073730469 + j-0.976989746094
            im_multiplicator=>-16007
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1101),
            data_im_in=>first_stage_im_out(1101),
            product_re_out=>mul_re_out(1101),
            product_im_out=>mul_im_out(1101)
        );

    UMUL_1102 : complex_multiplier
    generic map(
            re_multiplicator=>1805, --- 0.110168457031 + j-0.993896484375
            im_multiplicator=>-16284
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1102),
            data_im_in=>first_stage_im_out(1102),
            product_re_out=>mul_re_out(1102),
            product_im_out=>mul_im_out(1102)
        );

    UMUL_1103 : complex_multiplier
    generic map(
            re_multiplicator=>100, --- 0.006103515625 + j-0.999938964844
            im_multiplicator=>-16383
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1103),
            data_im_in=>first_stage_im_out(1103),
            product_re_out=>mul_re_out(1103),
            product_im_out=>mul_im_out(1103)
        );

    UMUL_1104 : complex_multiplier
    generic map(
            re_multiplicator=>-1605, --- -0.0979614257812 + j-0.995178222656
            im_multiplicator=>-16305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1104),
            data_im_in=>first_stage_im_out(1104),
            product_re_out=>mul_re_out(1104),
            product_im_out=>mul_im_out(1104)
        );

    UMUL_1105 : complex_multiplier
    generic map(
            re_multiplicator=>-3294, --- -0.201049804688 + j-0.979553222656
            im_multiplicator=>-16049
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1105),
            data_im_in=>first_stage_im_out(1105),
            product_re_out=>mul_re_out(1105),
            product_im_out=>mul_im_out(1105)
        );

    UMUL_1106 : complex_multiplier
    generic map(
            re_multiplicator=>-4948, --- -0.302001953125 + j-0.953247070312
            im_multiplicator=>-15618
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1106),
            data_im_in=>first_stage_im_out(1106),
            product_re_out=>mul_re_out(1106),
            product_im_out=>mul_im_out(1106)
        );

    UMUL_1107 : complex_multiplier
    generic map(
            re_multiplicator=>-6547, --- -0.399597167969 + j-0.916625976562
            im_multiplicator=>-15018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1107),
            data_im_in=>first_stage_im_out(1107),
            product_re_out=>mul_re_out(1107),
            product_im_out=>mul_im_out(1107)
        );

    UMUL_1108 : complex_multiplier
    generic map(
            re_multiplicator=>-8075, --- -0.492858886719 + j-0.870056152344
            im_multiplicator=>-14255
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1108),
            data_im_in=>first_stage_im_out(1108),
            product_re_out=>mul_re_out(1108),
            product_im_out=>mul_im_out(1108)
        );

    UMUL_1109 : complex_multiplier
    generic map(
            re_multiplicator=>-9516, --- -0.580810546875 + j-0.814025878906
            im_multiplicator=>-13337
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1109),
            data_im_in=>first_stage_im_out(1109),
            product_re_out=>mul_re_out(1109),
            product_im_out=>mul_im_out(1109)
        );

    UMUL_1110 : complex_multiplier
    generic map(
            re_multiplicator=>-10853, --- -0.662414550781 + j-0.749084472656
            im_multiplicator=>-12273
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1110),
            data_im_in=>first_stage_im_out(1110),
            product_re_out=>mul_re_out(1110),
            product_im_out=>mul_im_out(1110)
        );

    UMUL_1111 : complex_multiplier
    generic map(
            re_multiplicator=>-12072, --- -0.73681640625 + j-0.676086425781
            im_multiplicator=>-11077
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1111),
            data_im_in=>first_stage_im_out(1111),
            product_re_out=>mul_re_out(1111),
            product_im_out=>mul_im_out(1111)
        );

    UMUL_1112 : complex_multiplier
    generic map(
            re_multiplicator=>-13159, --- -0.803161621094 + j-0.595642089844
            im_multiplicator=>-9759
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1112),
            data_im_in=>first_stage_im_out(1112),
            product_re_out=>mul_re_out(1112),
            product_im_out=>mul_im_out(1112)
        );

    UMUL_1113 : complex_multiplier
    generic map(
            re_multiplicator=>-14104, --- -0.86083984375 + j-0.5087890625
            im_multiplicator=>-8336
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1113),
            data_im_in=>first_stage_im_out(1113),
            product_re_out=>mul_re_out(1113),
            product_im_out=>mul_im_out(1113)
        );

    UMUL_1114 : complex_multiplier
    generic map(
            re_multiplicator=>-14895, --- -0.909118652344 + j-0.416381835938
            im_multiplicator=>-6822
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1114),
            data_im_in=>first_stage_im_out(1114),
            product_re_out=>mul_re_out(1114),
            product_im_out=>mul_im_out(1114)
        );

    UMUL_1115 : complex_multiplier
    generic map(
            re_multiplicator=>-15525, --- -0.947570800781 + j-0.319458007812
            im_multiplicator=>-5234
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1115),
            data_im_in=>first_stage_im_out(1115),
            product_re_out=>mul_re_out(1115),
            product_im_out=>mul_im_out(1115)
        );

    UMUL_1116 : complex_multiplier
    generic map(
            re_multiplicator=>-15985, --- -0.975646972656 + j-0.219055175781
            im_multiplicator=>-3589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1116),
            data_im_in=>first_stage_im_out(1116),
            product_re_out=>mul_re_out(1116),
            product_im_out=>mul_im_out(1116)
        );

    UMUL_1117 : complex_multiplier
    generic map(
            re_multiplicator=>-16272, --- -0.9931640625 + j-0.116271972656
            im_multiplicator=>-1905
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1117),
            data_im_in=>first_stage_im_out(1117),
            product_re_out=>mul_re_out(1117),
            product_im_out=>mul_im_out(1117)
        );

    UMUL_1118 : complex_multiplier
    generic map(
            re_multiplicator=>-16382, --- -0.999877929688 + j-0.0122680664062
            im_multiplicator=>-201
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1118),
            data_im_in=>first_stage_im_out(1118),
            product_re_out=>mul_re_out(1118),
            product_im_out=>mul_im_out(1118)
        );

    UMUL_1119 : complex_multiplier
    generic map(
            re_multiplicator=>-16314, --- -0.995727539062 + j0.0918579101562
            im_multiplicator=>1505
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1119),
            data_im_in=>first_stage_im_out(1119),
            product_re_out=>mul_re_out(1119),
            product_im_out=>mul_im_out(1119)
        );

    UDELAY_1120_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1120),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1120)
        );
    UDELAY_1120_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1120),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1120)
        );
    USHIFTER_1120_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1120),
            data_out=>mul_re_out(1120)
        );
    USHIFTER_1120_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1120),
            data_out=>mul_im_out(1120)
        );

    UMUL_1121 : complex_multiplier
    generic map(
            re_multiplicator=>16289, --- 0.994201660156 + j-0.107116699219
            im_multiplicator=>-1755
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1121),
            data_im_in=>first_stage_im_out(1121),
            product_re_out=>mul_re_out(1121),
            product_im_out=>mul_im_out(1121)
        );

    UMUL_1122 : complex_multiplier
    generic map(
            re_multiplicator=>16007, --- 0.976989746094 + j-0.213073730469
            im_multiplicator=>-3491
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1122),
            data_im_in=>first_stage_im_out(1122),
            product_re_out=>mul_re_out(1122),
            product_im_out=>mul_im_out(1122)
        );

    UMUL_1123 : complex_multiplier
    generic map(
            re_multiplicator=>15541, --- 0.948547363281 + j-0.316589355469
            im_multiplicator=>-5187
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1123),
            data_im_in=>first_stage_im_out(1123),
            product_re_out=>mul_re_out(1123),
            product_im_out=>mul_im_out(1123)
        );

    UMUL_1124 : complex_multiplier
    generic map(
            re_multiplicator=>14895, --- 0.909118652344 + j-0.416381835938
            im_multiplicator=>-6822
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1124),
            data_im_in=>first_stage_im_out(1124),
            product_re_out=>mul_re_out(1124),
            product_im_out=>mul_im_out(1124)
        );

    UMUL_1125 : complex_multiplier
    generic map(
            re_multiplicator=>14078, --- 0.859252929688 + j-0.511413574219
            im_multiplicator=>-8379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1125),
            data_im_in=>first_stage_im_out(1125),
            product_re_out=>mul_re_out(1125),
            product_im_out=>mul_im_out(1125)
        );

    UMUL_1126 : complex_multiplier
    generic map(
            re_multiplicator=>13099, --- 0.799499511719 + j-0.6005859375
            im_multiplicator=>-9840
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1126),
            data_im_in=>first_stage_im_out(1126),
            product_re_out=>mul_re_out(1126),
            product_im_out=>mul_im_out(1126)
        );

    UMUL_1127 : complex_multiplier
    generic map(
            re_multiplicator=>11969, --- 0.730529785156 + j-0.682800292969
            im_multiplicator=>-11187
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1127),
            data_im_in=>first_stage_im_out(1127),
            product_re_out=>mul_re_out(1127),
            product_im_out=>mul_im_out(1127)
        );

    UMUL_1128 : complex_multiplier
    generic map(
            re_multiplicator=>10701, --- 0.653137207031 + j-0.757202148438
            im_multiplicator=>-12406
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1128),
            data_im_in=>first_stage_im_out(1128),
            product_re_out=>mul_re_out(1128),
            product_im_out=>mul_im_out(1128)
        );

    UMUL_1129 : complex_multiplier
    generic map(
            re_multiplicator=>9310, --- 0.568237304688 + j-0.822814941406
            im_multiplicator=>-13481
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1129),
            data_im_in=>first_stage_im_out(1129),
            product_re_out=>mul_re_out(1129),
            product_im_out=>mul_im_out(1129)
        );

    UMUL_1130 : complex_multiplier
    generic map(
            re_multiplicator=>7811, --- 0.476745605469 + j-0.878967285156
            im_multiplicator=>-14401
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1130),
            data_im_in=>first_stage_im_out(1130),
            product_re_out=>mul_re_out(1130),
            product_im_out=>mul_im_out(1130)
        );

    UMUL_1131 : complex_multiplier
    generic map(
            re_multiplicator=>6223, --- 0.379821777344 + j-0.925048828125
            im_multiplicator=>-15156
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1131),
            data_im_in=>first_stage_im_out(1131),
            product_re_out=>mul_re_out(1131),
            product_im_out=>mul_im_out(1131)
        );

    UMUL_1132 : complex_multiplier
    generic map(
            re_multiplicator=>4563, --- 0.278503417969 + j-0.960388183594
            im_multiplicator=>-15735
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1132),
            data_im_in=>first_stage_im_out(1132),
            product_re_out=>mul_re_out(1132),
            product_im_out=>mul_im_out(1132)
        );

    UMUL_1133 : complex_multiplier
    generic map(
            re_multiplicator=>2850, --- 0.173950195312 + j-0.984741210938
            im_multiplicator=>-16134
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1133),
            data_im_in=>first_stage_im_out(1133),
            product_re_out=>mul_re_out(1133),
            product_im_out=>mul_im_out(1133)
        );

    UMUL_1134 : complex_multiplier
    generic map(
            re_multiplicator=>1105, --- 0.0674438476562 + j-0.997680664062
            im_multiplicator=>-16346
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1134),
            data_im_in=>first_stage_im_out(1134),
            product_re_out=>mul_re_out(1134),
            product_im_out=>mul_im_out(1134)
        );

    UMUL_1135 : complex_multiplier
    generic map(
            re_multiplicator=>-653, --- -0.0398559570312 + j-0.999145507812
            im_multiplicator=>-16370
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1135),
            data_im_in=>first_stage_im_out(1135),
            product_re_out=>mul_re_out(1135),
            product_im_out=>mul_im_out(1135)
        );

    UMUL_1136 : complex_multiplier
    generic map(
            re_multiplicator=>-2404, --- -0.146728515625 + j-0.989135742188
            im_multiplicator=>-16206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1136),
            data_im_in=>first_stage_im_out(1136),
            product_re_out=>mul_re_out(1136),
            product_im_out=>mul_im_out(1136)
        );

    UMUL_1137 : complex_multiplier
    generic map(
            re_multiplicator=>-4127, --- -0.251892089844 + j-0.967712402344
            im_multiplicator=>-15855
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1137),
            data_im_in=>first_stage_im_out(1137),
            product_re_out=>mul_re_out(1137),
            product_im_out=>mul_im_out(1137)
        );

    UMUL_1138 : complex_multiplier
    generic map(
            re_multiplicator=>-5802, --- -0.354125976562 + j-0.935180664062
            im_multiplicator=>-15322
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1138),
            data_im_in=>first_stage_im_out(1138),
            product_re_out=>mul_re_out(1138),
            product_im_out=>mul_im_out(1138)
        );

    UMUL_1139 : complex_multiplier
    generic map(
            re_multiplicator=>-7411, --- -0.452331542969 + j-0.891784667969
            im_multiplicator=>-14611
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1139),
            data_im_in=>first_stage_im_out(1139),
            product_re_out=>mul_re_out(1139),
            product_im_out=>mul_im_out(1139)
        );

    UMUL_1140 : complex_multiplier
    generic map(
            re_multiplicator=>-8934, --- -0.545288085938 + j-0.838195800781
            im_multiplicator=>-13733
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1140),
            data_im_in=>first_stage_im_out(1140),
            product_re_out=>mul_re_out(1140),
            product_im_out=>mul_im_out(1140)
        );

    UMUL_1141 : complex_multiplier
    generic map(
            re_multiplicator=>-10354, --- -0.631958007812 + j-0.77490234375
            im_multiplicator=>-12696
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1141),
            data_im_in=>first_stage_im_out(1141),
            product_re_out=>mul_re_out(1141),
            product_im_out=>mul_im_out(1141)
        );

    UMUL_1142 : complex_multiplier
    generic map(
            re_multiplicator=>-11656, --- -0.71142578125 + j-0.702697753906
            im_multiplicator=>-11513
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1142),
            data_im_in=>first_stage_im_out(1142),
            product_re_out=>mul_re_out(1142),
            product_im_out=>mul_im_out(1142)
        );

    UMUL_1143 : complex_multiplier
    generic map(
            re_multiplicator=>-12822, --- -0.782592773438 + j-0.622436523438
            im_multiplicator=>-10198
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1143),
            data_im_in=>first_stage_im_out(1143),
            product_re_out=>mul_re_out(1143),
            product_im_out=>mul_im_out(1143)
        );

    UMUL_1144 : complex_multiplier
    generic map(
            re_multiplicator=>-13842, --- -0.844848632812 + j-0.534973144531
            im_multiplicator=>-8765
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1144),
            data_im_in=>first_stage_im_out(1144),
            product_re_out=>mul_re_out(1144),
            product_im_out=>mul_im_out(1144)
        );

    UMUL_1145 : complex_multiplier
    generic map(
            re_multiplicator=>-14701, --- -0.897277832031 + j-0.441345214844
            im_multiplicator=>-7231
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1145),
            data_im_in=>first_stage_im_out(1145),
            product_re_out=>mul_re_out(1145),
            product_im_out=>mul_im_out(1145)
        );

    UMUL_1146 : complex_multiplier
    generic map(
            re_multiplicator=>-15392, --- -0.939453125 + j-0.342651367188
            im_multiplicator=>-5614
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1146),
            data_im_in=>first_stage_im_out(1146),
            product_re_out=>mul_re_out(1146),
            product_im_out=>mul_im_out(1146)
        );

    UMUL_1147 : complex_multiplier
    generic map(
            re_multiplicator=>-15905, --- -0.970764160156 + j-0.239990234375
            im_multiplicator=>-3932
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1147),
            data_im_in=>first_stage_im_out(1147),
            product_re_out=>mul_re_out(1147),
            product_im_out=>mul_im_out(1147)
        );

    UMUL_1148 : complex_multiplier
    generic map(
            re_multiplicator=>-16234, --- -0.990844726562 + j-0.134521484375
            im_multiplicator=>-2204
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1148),
            data_im_in=>first_stage_im_out(1148),
            product_re_out=>mul_re_out(1148),
            product_im_out=>mul_im_out(1148)
        );

    UMUL_1149 : complex_multiplier
    generic map(
            re_multiplicator=>-16377, --- -0.999572753906 + j-0.027587890625
            im_multiplicator=>-452
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1149),
            data_im_in=>first_stage_im_out(1149),
            product_re_out=>mul_re_out(1149),
            product_im_out=>mul_im_out(1149)
        );

    UMUL_1150 : complex_multiplier
    generic map(
            re_multiplicator=>-16331, --- -0.996765136719 + j0.0796508789062
            im_multiplicator=>1305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1150),
            data_im_in=>first_stage_im_out(1150),
            product_re_out=>mul_re_out(1150),
            product_im_out=>mul_im_out(1150)
        );

    UMUL_1151 : complex_multiplier
    generic map(
            re_multiplicator=>-16097, --- -0.982482910156 + j0.18603515625
            im_multiplicator=>3048
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1151),
            data_im_in=>first_stage_im_out(1151),
            product_re_out=>mul_re_out(1151),
            product_im_out=>mul_im_out(1151)
        );

    UDELAY_1152_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1152),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1152)
        );
    UDELAY_1152_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1152),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1152)
        );
    USHIFTER_1152_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1152),
            data_out=>mul_re_out(1152)
        );
    USHIFTER_1152_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1152),
            data_out=>mul_im_out(1152)
        );

    UMUL_1153 : complex_multiplier
    generic map(
            re_multiplicator=>16284, --- 0.993896484375 + j-0.110168457031
            im_multiplicator=>-1805
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1153),
            data_im_in=>first_stage_im_out(1153),
            product_re_out=>mul_re_out(1153),
            product_im_out=>mul_im_out(1153)
        );

    UMUL_1154 : complex_multiplier
    generic map(
            re_multiplicator=>15985, --- 0.975646972656 + j-0.219055175781
            im_multiplicator=>-3589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1154),
            data_im_in=>first_stage_im_out(1154),
            product_re_out=>mul_re_out(1154),
            product_im_out=>mul_im_out(1154)
        );

    UMUL_1155 : complex_multiplier
    generic map(
            re_multiplicator=>15492, --- 0.945556640625 + j-0.325256347656
            im_multiplicator=>-5329
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1155),
            data_im_in=>first_stage_im_out(1155),
            product_re_out=>mul_re_out(1155),
            product_im_out=>mul_im_out(1155)
        );

    UMUL_1156 : complex_multiplier
    generic map(
            re_multiplicator=>14810, --- 0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1156),
            data_im_in=>first_stage_im_out(1156),
            product_re_out=>mul_re_out(1156),
            product_im_out=>mul_im_out(1156)
        );

    UMUL_1157 : complex_multiplier
    generic map(
            re_multiplicator=>13948, --- 0.851318359375 + j-0.524536132812
            im_multiplicator=>-8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1157),
            data_im_in=>first_stage_im_out(1157),
            product_re_out=>mul_re_out(1157),
            product_im_out=>mul_im_out(1157)
        );

    UMUL_1158 : complex_multiplier
    generic map(
            re_multiplicator=>12916, --- 0.788330078125 + j-0.615173339844
            im_multiplicator=>-10079
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1158),
            data_im_in=>first_stage_im_out(1158),
            product_re_out=>mul_re_out(1158),
            product_im_out=>mul_im_out(1158)
        );

    UMUL_1159 : complex_multiplier
    generic map(
            re_multiplicator=>11726, --- 0.715698242188 + j-0.698364257812
            im_multiplicator=>-11442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1159),
            data_im_in=>first_stage_im_out(1159),
            product_re_out=>mul_re_out(1159),
            product_im_out=>mul_im_out(1159)
        );

    UMUL_1160 : complex_multiplier
    generic map(
            re_multiplicator=>10393, --- 0.634338378906 + j-0.773010253906
            im_multiplicator=>-12665
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1160),
            data_im_in=>first_stage_im_out(1160),
            product_re_out=>mul_re_out(1160),
            product_im_out=>mul_im_out(1160)
        );

    UMUL_1161 : complex_multiplier
    generic map(
            re_multiplicator=>8934, --- 0.545288085938 + j-0.838195800781
            im_multiplicator=>-13733
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1161),
            data_im_in=>first_stage_im_out(1161),
            product_re_out=>mul_re_out(1161),
            product_im_out=>mul_im_out(1161)
        );

    UMUL_1162 : complex_multiplier
    generic map(
            re_multiplicator=>7366, --- 0.449584960938 + j-0.893188476562
            im_multiplicator=>-14634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1162),
            data_im_in=>first_stage_im_out(1162),
            product_re_out=>mul_re_out(1162),
            product_im_out=>mul_im_out(1162)
        );

    UMUL_1163 : complex_multiplier
    generic map(
            re_multiplicator=>5708, --- 0.348388671875 + j-0.937316894531
            im_multiplicator=>-15357
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1163),
            data_im_in=>first_stage_im_out(1163),
            product_re_out=>mul_re_out(1163),
            product_im_out=>mul_im_out(1163)
        );

    UMUL_1164 : complex_multiplier
    generic map(
            re_multiplicator=>3980, --- 0.242919921875 + j-0.969970703125
            im_multiplicator=>-15892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1164),
            data_im_in=>first_stage_im_out(1164),
            product_re_out=>mul_re_out(1164),
            product_im_out=>mul_im_out(1164)
        );

    UMUL_1165 : complex_multiplier
    generic map(
            re_multiplicator=>2204, --- 0.134521484375 + j-0.990844726562
            im_multiplicator=>-16234
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1165),
            data_im_in=>first_stage_im_out(1165),
            product_re_out=>mul_re_out(1165),
            product_im_out=>mul_im_out(1165)
        );

    UMUL_1166 : complex_multiplier
    generic map(
            re_multiplicator=>402, --- 0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1166),
            data_im_in=>first_stage_im_out(1166),
            product_re_out=>mul_re_out(1166),
            product_im_out=>mul_im_out(1166)
        );

    UMUL_1167 : complex_multiplier
    generic map(
            re_multiplicator=>-1405, --- -0.0857543945312 + j-0.996276855469
            im_multiplicator=>-16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1167),
            data_im_in=>first_stage_im_out(1167),
            product_re_out=>mul_re_out(1167),
            product_im_out=>mul_im_out(1167)
        );

    UMUL_1168 : complex_multiplier
    generic map(
            re_multiplicator=>-3196, --- -0.195068359375 + j-0.980773925781
            im_multiplicator=>-16069
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1168),
            data_im_in=>first_stage_im_out(1168),
            product_re_out=>mul_re_out(1168),
            product_im_out=>mul_im_out(1168)
        );

    UMUL_1169 : complex_multiplier
    generic map(
            re_multiplicator=>-4948, --- -0.302001953125 + j-0.953247070312
            im_multiplicator=>-15618
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1169),
            data_im_in=>first_stage_im_out(1169),
            product_re_out=>mul_re_out(1169),
            product_im_out=>mul_im_out(1169)
        );

    UMUL_1170 : complex_multiplier
    generic map(
            re_multiplicator=>-6639, --- -0.405212402344 + j-0.914184570312
            im_multiplicator=>-14978
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1170),
            data_im_in=>first_stage_im_out(1170),
            product_re_out=>mul_re_out(1170),
            product_im_out=>mul_im_out(1170)
        );

    UMUL_1171 : complex_multiplier
    generic map(
            re_multiplicator=>-8249, --- -0.503479003906 + j-0.863952636719
            im_multiplicator=>-14155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1171),
            data_im_in=>first_stage_im_out(1171),
            product_re_out=>mul_re_out(1171),
            product_im_out=>mul_im_out(1171)
        );

    UMUL_1172 : complex_multiplier
    generic map(
            re_multiplicator=>-9759, --- -0.595642089844 + j-0.803161621094
            im_multiplicator=>-13159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1172),
            data_im_in=>first_stage_im_out(1172),
            product_re_out=>mul_re_out(1172),
            product_im_out=>mul_im_out(1172)
        );

    UMUL_1173 : complex_multiplier
    generic map(
            re_multiplicator=>-11150, --- -0.680541992188 + j-0.732604980469
            im_multiplicator=>-12003
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1173),
            data_im_in=>first_stage_im_out(1173),
            product_re_out=>mul_re_out(1173),
            product_im_out=>mul_im_out(1173)
        );

    UMUL_1174 : complex_multiplier
    generic map(
            re_multiplicator=>-12406, --- -0.757202148438 + j-0.653137207031
            im_multiplicator=>-10701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1174),
            data_im_in=>first_stage_im_out(1174),
            product_re_out=>mul_re_out(1174),
            product_im_out=>mul_im_out(1174)
        );

    UMUL_1175 : complex_multiplier
    generic map(
            re_multiplicator=>-13510, --- -0.824584960938 + j-0.565673828125
            im_multiplicator=>-9268
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1175),
            data_im_in=>first_stage_im_out(1175),
            product_re_out=>mul_re_out(1175),
            product_im_out=>mul_im_out(1175)
        );

    UMUL_1176 : complex_multiplier
    generic map(
            re_multiplicator=>-14449, --- -0.881896972656 + j-0.471374511719
            im_multiplicator=>-7723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1176),
            data_im_in=>first_stage_im_out(1176),
            product_re_out=>mul_re_out(1176),
            product_im_out=>mul_im_out(1176)
        );

    UMUL_1177 : complex_multiplier
    generic map(
            re_multiplicator=>-15212, --- -0.928466796875 + j-0.371276855469
            im_multiplicator=>-6083
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1177),
            data_im_in=>first_stage_im_out(1177),
            product_re_out=>mul_re_out(1177),
            product_im_out=>mul_im_out(1177)
        );

    UMUL_1178 : complex_multiplier
    generic map(
            re_multiplicator=>-15790, --- -0.963745117188 + j-0.266662597656
            im_multiplicator=>-4369
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1178),
            data_im_in=>first_stage_im_out(1178),
            product_re_out=>mul_re_out(1178),
            product_im_out=>mul_im_out(1178)
        );

    UMUL_1179 : complex_multiplier
    generic map(
            re_multiplicator=>-16175, --- -0.987243652344 + j-0.158813476562
            im_multiplicator=>-2602
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1179),
            data_im_in=>first_stage_im_out(1179),
            product_re_out=>mul_re_out(1179),
            product_im_out=>mul_im_out(1179)
        );

    UMUL_1180 : complex_multiplier
    generic map(
            re_multiplicator=>-16364, --- -0.998779296875 + j-0.0490112304688
            im_multiplicator=>-803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1180),
            data_im_in=>first_stage_im_out(1180),
            product_re_out=>mul_re_out(1180),
            product_im_out=>mul_im_out(1180)
        );

    UMUL_1181 : complex_multiplier
    generic map(
            re_multiplicator=>-16353, --- -0.998107910156 + j0.061279296875
            im_multiplicator=>1004
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1181),
            data_im_in=>first_stage_im_out(1181),
            product_re_out=>mul_re_out(1181),
            product_im_out=>mul_im_out(1181)
        );

    UMUL_1182 : complex_multiplier
    generic map(
            re_multiplicator=>-16142, --- -0.985229492188 + j0.170959472656
            im_multiplicator=>2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1182),
            data_im_in=>first_stage_im_out(1182),
            product_re_out=>mul_re_out(1182),
            product_im_out=>mul_im_out(1182)
        );

    UMUL_1183 : complex_multiplier
    generic map(
            re_multiplicator=>-15735, --- -0.960388183594 + j0.278503417969
            im_multiplicator=>4563
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1183),
            data_im_in=>first_stage_im_out(1183),
            product_re_out=>mul_re_out(1183),
            product_im_out=>mul_im_out(1183)
        );

    UDELAY_1184_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1184),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1184)
        );
    UDELAY_1184_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1184),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1184)
        );
    USHIFTER_1184_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1184),
            data_out=>mul_re_out(1184)
        );
    USHIFTER_1184_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1184),
            data_out=>mul_im_out(1184)
        );

    UMUL_1185 : complex_multiplier
    generic map(
            re_multiplicator=>16278, --- 0.993530273438 + j-0.113220214844
            im_multiplicator=>-1855
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1185),
            data_im_in=>first_stage_im_out(1185),
            product_re_out=>mul_re_out(1185),
            product_im_out=>mul_im_out(1185)
        );

    UMUL_1186 : complex_multiplier
    generic map(
            re_multiplicator=>15963, --- 0.974304199219 + j-0.225036621094
            im_multiplicator=>-3687
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1186),
            data_im_in=>first_stage_im_out(1186),
            product_re_out=>mul_re_out(1186),
            product_im_out=>mul_im_out(1186)
        );

    UMUL_1187 : complex_multiplier
    generic map(
            re_multiplicator=>15443, --- 0.942565917969 + j-0.333984375
            im_multiplicator=>-5472
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1187),
            data_im_in=>first_stage_im_out(1187),
            product_re_out=>mul_re_out(1187),
            product_im_out=>mul_im_out(1187)
        );

    UMUL_1188 : complex_multiplier
    generic map(
            re_multiplicator=>14723, --- 0.898620605469 + j-0.438598632812
            im_multiplicator=>-7186
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1188),
            data_im_in=>first_stage_im_out(1188),
            product_re_out=>mul_re_out(1188),
            product_im_out=>mul_im_out(1188)
        );

    UMUL_1189 : complex_multiplier
    generic map(
            re_multiplicator=>13815, --- 0.843200683594 + j-0.537536621094
            im_multiplicator=>-8807
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1189),
            data_im_in=>first_stage_im_out(1189),
            product_re_out=>mul_re_out(1189),
            product_im_out=>mul_im_out(1189)
        );

    UMUL_1190 : complex_multiplier
    generic map(
            re_multiplicator=>12728, --- 0.77685546875 + j-0.629577636719
            im_multiplicator=>-10315
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1190),
            data_im_in=>first_stage_im_out(1190),
            product_re_out=>mul_re_out(1190),
            product_im_out=>mul_im_out(1190)
        );

    UMUL_1191 : complex_multiplier
    generic map(
            re_multiplicator=>11478, --- 0.700561523438 + j-0.713562011719
            im_multiplicator=>-11691
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1191),
            data_im_in=>first_stage_im_out(1191),
            product_re_out=>mul_re_out(1191),
            product_im_out=>mul_im_out(1191)
        );

    UMUL_1192 : complex_multiplier
    generic map(
            re_multiplicator=>10079, --- 0.615173339844 + j-0.788330078125
            im_multiplicator=>-12916
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1192),
            data_im_in=>first_stage_im_out(1192),
            product_re_out=>mul_re_out(1192),
            product_im_out=>mul_im_out(1192)
        );

    UMUL_1193 : complex_multiplier
    generic map(
            re_multiplicator=>8552, --- 0.52197265625 + j-0.852905273438
            im_multiplicator=>-13974
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1193),
            data_im_in=>first_stage_im_out(1193),
            product_re_out=>mul_re_out(1193),
            product_im_out=>mul_im_out(1193)
        );

    UMUL_1194 : complex_multiplier
    generic map(
            re_multiplicator=>6914, --- 0.421997070312 + j-0.906555175781
            im_multiplicator=>-14853
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1194),
            data_im_in=>first_stage_im_out(1194),
            product_re_out=>mul_re_out(1194),
            product_im_out=>mul_im_out(1194)
        );

    UMUL_1195 : complex_multiplier
    generic map(
            re_multiplicator=>5187, --- 0.316589355469 + j-0.948547363281
            im_multiplicator=>-15541
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1195),
            data_im_in=>first_stage_im_out(1195),
            product_re_out=>mul_re_out(1195),
            product_im_out=>mul_im_out(1195)
        );

    UMUL_1196 : complex_multiplier
    generic map(
            re_multiplicator=>3393, --- 0.207092285156 + j-0.978271484375
            im_multiplicator=>-16028
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1196),
            data_im_in=>first_stage_im_out(1196),
            product_re_out=>mul_re_out(1196),
            product_im_out=>mul_im_out(1196)
        );

    UMUL_1197 : complex_multiplier
    generic map(
            re_multiplicator=>1555, --- 0.0949096679688 + j-0.995422363281
            im_multiplicator=>-16309
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1197),
            data_im_in=>first_stage_im_out(1197),
            product_re_out=>mul_re_out(1197),
            product_im_out=>mul_im_out(1197)
        );

    UMUL_1198 : complex_multiplier
    generic map(
            re_multiplicator=>-301, --- -0.0183715820312 + j-0.999816894531
            im_multiplicator=>-16381
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1198),
            data_im_in=>first_stage_im_out(1198),
            product_re_out=>mul_re_out(1198),
            product_im_out=>mul_im_out(1198)
        );

    UMUL_1199 : complex_multiplier
    generic map(
            re_multiplicator=>-2155, --- -0.131530761719 + j-0.991271972656
            im_multiplicator=>-16241
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1199),
            data_im_in=>first_stage_im_out(1199),
            product_re_out=>mul_re_out(1199),
            product_im_out=>mul_im_out(1199)
        );

    UMUL_1200 : complex_multiplier
    generic map(
            re_multiplicator=>-3980, --- -0.242919921875 + j-0.969970703125
            im_multiplicator=>-15892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1200),
            data_im_in=>first_stage_im_out(1200),
            product_re_out=>mul_re_out(1200),
            product_im_out=>mul_im_out(1200)
        );

    UMUL_1201 : complex_multiplier
    generic map(
            re_multiplicator=>-5755, --- -0.351257324219 + j-0.936218261719
            im_multiplicator=>-15339
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1201),
            data_im_in=>first_stage_im_out(1201),
            product_re_out=>mul_re_out(1201),
            product_im_out=>mul_im_out(1201)
        );

    UMUL_1202 : complex_multiplier
    generic map(
            re_multiplicator=>-7456, --- -0.455078125 + j-0.890441894531
            im_multiplicator=>-14589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1202),
            data_im_in=>first_stage_im_out(1202),
            product_re_out=>mul_re_out(1202),
            product_im_out=>mul_im_out(1202)
        );

    UMUL_1203 : complex_multiplier
    generic map(
            re_multiplicator=>-9060, --- -0.552978515625 + j-0.833129882812
            im_multiplicator=>-13650
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1203),
            data_im_in=>first_stage_im_out(1203),
            product_re_out=>mul_re_out(1203),
            product_im_out=>mul_im_out(1203)
        );

    UMUL_1204 : complex_multiplier
    generic map(
            re_multiplicator=>-10548, --- -0.643798828125 + j-0.76513671875
            im_multiplicator=>-12536
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1204),
            data_im_in=>first_stage_im_out(1204),
            product_re_out=>mul_re_out(1204),
            product_im_out=>mul_im_out(1204)
        );

    UMUL_1205 : complex_multiplier
    generic map(
            re_multiplicator=>-11900, --- -0.726318359375 + j-0.687255859375
            im_multiplicator=>-11260
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1205),
            data_im_in=>first_stage_im_out(1205),
            product_re_out=>mul_re_out(1205),
            product_im_out=>mul_im_out(1205)
        );

    UMUL_1206 : complex_multiplier
    generic map(
            re_multiplicator=>-13099, --- -0.799499511719 + j-0.6005859375
            im_multiplicator=>-9840
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1206),
            data_im_in=>first_stage_im_out(1206),
            product_re_out=>mul_re_out(1206),
            product_im_out=>mul_im_out(1206)
        );

    UMUL_1207 : complex_multiplier
    generic map(
            re_multiplicator=>-14129, --- -0.862365722656 + j-0.506164550781
            im_multiplicator=>-8293
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1207),
            data_im_in=>first_stage_im_out(1207),
            product_re_out=>mul_re_out(1207),
            product_im_out=>mul_im_out(1207)
        );

    UMUL_1208 : complex_multiplier
    generic map(
            re_multiplicator=>-14978, --- -0.914184570312 + j-0.405212402344
            im_multiplicator=>-6639
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1208),
            data_im_in=>first_stage_im_out(1208),
            product_re_out=>mul_re_out(1208),
            product_im_out=>mul_im_out(1208)
        );

    UMUL_1209 : complex_multiplier
    generic map(
            re_multiplicator=>-15634, --- -0.954223632812 + j-0.299072265625
            im_multiplicator=>-4900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1209),
            data_im_in=>first_stage_im_out(1209),
            product_re_out=>mul_re_out(1209),
            product_im_out=>mul_im_out(1209)
        );

    UMUL_1210 : complex_multiplier
    generic map(
            re_multiplicator=>-16088, --- -0.98193359375 + j-0.189025878906
            im_multiplicator=>-3097
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1210),
            data_im_in=>first_stage_im_out(1210),
            product_re_out=>mul_re_out(1210),
            product_im_out=>mul_im_out(1210)
        );

    UMUL_1211 : complex_multiplier
    generic map(
            re_multiplicator=>-16335, --- -0.997009277344 + j-0.0765991210938
            im_multiplicator=>-1255
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1211),
            data_im_in=>first_stage_im_out(1211),
            product_re_out=>mul_re_out(1211),
            product_im_out=>mul_im_out(1211)
        );

    UMUL_1212 : complex_multiplier
    generic map(
            re_multiplicator=>-16372, --- -0.999267578125 + j0.0368041992188
            im_multiplicator=>603
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1212),
            data_im_in=>first_stage_im_out(1212),
            product_re_out=>mul_re_out(1212),
            product_im_out=>mul_im_out(1212)
        );

    UMUL_1213 : complex_multiplier
    generic map(
            re_multiplicator=>-16199, --- -0.988708496094 + j0.149719238281
            im_multiplicator=>2453
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1213),
            data_im_in=>first_stage_im_out(1213),
            product_re_out=>mul_re_out(1213),
            product_im_out=>mul_im_out(1213)
        );

    UMUL_1214 : complex_multiplier
    generic map(
            re_multiplicator=>-15817, --- -0.965393066406 + j0.2607421875
            im_multiplicator=>4272
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1214),
            data_im_in=>first_stage_im_out(1214),
            product_re_out=>mul_re_out(1214),
            product_im_out=>mul_im_out(1214)
        );

    UMUL_1215 : complex_multiplier
    generic map(
            re_multiplicator=>-15231, --- -0.929626464844 + j0.368408203125
            im_multiplicator=>6036
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1215),
            data_im_in=>first_stage_im_out(1215),
            product_re_out=>mul_re_out(1215),
            product_im_out=>mul_im_out(1215)
        );

    UDELAY_1216_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1216),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1216)
        );
    UDELAY_1216_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1216),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1216)
        );
    USHIFTER_1216_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1216),
            data_out=>mul_re_out(1216)
        );
    USHIFTER_1216_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1216),
            data_out=>mul_im_out(1216)
        );

    UMUL_1217 : complex_multiplier
    generic map(
            re_multiplicator=>16272, --- 0.9931640625 + j-0.116271972656
            im_multiplicator=>-1905
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1217),
            data_im_in=>first_stage_im_out(1217),
            product_re_out=>mul_re_out(1217),
            product_im_out=>mul_im_out(1217)
        );

    UMUL_1218 : complex_multiplier
    generic map(
            re_multiplicator=>15940, --- 0.972900390625 + j-0.231018066406
            im_multiplicator=>-3785
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1218),
            data_im_in=>first_stage_im_out(1218),
            product_re_out=>mul_re_out(1218),
            product_im_out=>mul_im_out(1218)
        );

    UMUL_1219 : complex_multiplier
    generic map(
            re_multiplicator=>15392, --- 0.939453125 + j-0.342651367188
            im_multiplicator=>-5614
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1219),
            data_im_in=>first_stage_im_out(1219),
            product_re_out=>mul_re_out(1219),
            product_im_out=>mul_im_out(1219)
        );

    UMUL_1220 : complex_multiplier
    generic map(
            re_multiplicator=>14634, --- 0.893188476562 + j-0.449584960938
            im_multiplicator=>-7366
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1220),
            data_im_in=>first_stage_im_out(1220),
            product_re_out=>mul_re_out(1220),
            product_im_out=>mul_im_out(1220)
        );

    UMUL_1221 : complex_multiplier
    generic map(
            re_multiplicator=>13678, --- 0.834838867188 + j-0.550415039062
            im_multiplicator=>-9018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1221),
            data_im_in=>first_stage_im_out(1221),
            product_re_out=>mul_re_out(1221),
            product_im_out=>mul_im_out(1221)
        );

    UMUL_1222 : complex_multiplier
    generic map(
            re_multiplicator=>12536, --- 0.76513671875 + j-0.643798828125
            im_multiplicator=>-10548
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1222),
            data_im_in=>first_stage_im_out(1222),
            product_re_out=>mul_re_out(1222),
            product_im_out=>mul_im_out(1222)
        );

    UMUL_1223 : complex_multiplier
    generic map(
            re_multiplicator=>11224, --- 0.68505859375 + j-0.728454589844
            im_multiplicator=>-11935
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1223),
            data_im_in=>first_stage_im_out(1223),
            product_re_out=>mul_re_out(1223),
            product_im_out=>mul_im_out(1223)
        );

    UMUL_1224 : complex_multiplier
    generic map(
            re_multiplicator=>9759, --- 0.595642089844 + j-0.803161621094
            im_multiplicator=>-13159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1224),
            data_im_in=>first_stage_im_out(1224),
            product_re_out=>mul_re_out(1224),
            product_im_out=>mul_im_out(1224)
        );

    UMUL_1225 : complex_multiplier
    generic map(
            re_multiplicator=>8162, --- 0.498168945312 + j-0.867004394531
            im_multiplicator=>-14205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1225),
            data_im_in=>first_stage_im_out(1225),
            product_re_out=>mul_re_out(1225),
            product_im_out=>mul_im_out(1225)
        );

    UMUL_1226 : complex_multiplier
    generic map(
            re_multiplicator=>6455, --- 0.393981933594 + j-0.919067382812
            im_multiplicator=>-15058
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1226),
            data_im_in=>first_stage_im_out(1226),
            product_re_out=>mul_re_out(1226),
            product_im_out=>mul_im_out(1226)
        );

    UMUL_1227 : complex_multiplier
    generic map(
            re_multiplicator=>4659, --- 0.284362792969 + j-0.958679199219
            im_multiplicator=>-15707
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1227),
            data_im_in=>first_stage_im_out(1227),
            product_re_out=>mul_re_out(1227),
            product_im_out=>mul_im_out(1227)
        );

    UMUL_1228 : complex_multiplier
    generic map(
            re_multiplicator=>2801, --- 0.170959472656 + j-0.985229492188
            im_multiplicator=>-16142
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1228),
            data_im_in=>first_stage_im_out(1228),
            product_re_out=>mul_re_out(1228),
            product_im_out=>mul_im_out(1228)
        );

    UMUL_1229 : complex_multiplier
    generic map(
            re_multiplicator=>904, --- 0.05517578125 + j-0.998474121094
            im_multiplicator=>-16359
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1229),
            data_im_in=>first_stage_im_out(1229),
            product_re_out=>mul_re_out(1229),
            product_im_out=>mul_im_out(1229)
        );

    UMUL_1230 : complex_multiplier
    generic map(
            re_multiplicator=>-1004, --- -0.061279296875 + j-0.998107910156
            im_multiplicator=>-16353
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1230),
            data_im_in=>first_stage_im_out(1230),
            product_re_out=>mul_re_out(1230),
            product_im_out=>mul_im_out(1230)
        );

    UMUL_1231 : complex_multiplier
    generic map(
            re_multiplicator=>-2900, --- -0.177001953125 + j-0.984191894531
            im_multiplicator=>-16125
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1231),
            data_im_in=>first_stage_im_out(1231),
            product_re_out=>mul_re_out(1231),
            product_im_out=>mul_im_out(1231)
        );

    UMUL_1232 : complex_multiplier
    generic map(
            re_multiplicator=>-4756, --- -0.290283203125 + j-0.956909179688
            im_multiplicator=>-15678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1232),
            data_im_in=>first_stage_im_out(1232),
            product_re_out=>mul_re_out(1232),
            product_im_out=>mul_im_out(1232)
        );

    UMUL_1233 : complex_multiplier
    generic map(
            re_multiplicator=>-6547, --- -0.399597167969 + j-0.916625976562
            im_multiplicator=>-15018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1233),
            data_im_in=>first_stage_im_out(1233),
            product_re_out=>mul_re_out(1233),
            product_im_out=>mul_im_out(1233)
        );

    UMUL_1234 : complex_multiplier
    generic map(
            re_multiplicator=>-8249, --- -0.503479003906 + j-0.863952636719
            im_multiplicator=>-14155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1234),
            data_im_in=>first_stage_im_out(1234),
            product_re_out=>mul_re_out(1234),
            product_im_out=>mul_im_out(1234)
        );

    UMUL_1235 : complex_multiplier
    generic map(
            re_multiplicator=>-9840, --- -0.6005859375 + j-0.799499511719
            im_multiplicator=>-13099
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1235),
            data_im_in=>first_stage_im_out(1235),
            product_re_out=>mul_re_out(1235),
            product_im_out=>mul_im_out(1235)
        );

    UMUL_1236 : complex_multiplier
    generic map(
            re_multiplicator=>-11297, --- -0.689514160156 + j-0.724243164062
            im_multiplicator=>-11866
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1236),
            data_im_in=>first_stage_im_out(1236),
            product_re_out=>mul_re_out(1236),
            product_im_out=>mul_im_out(1236)
        );

    UMUL_1237 : complex_multiplier
    generic map(
            re_multiplicator=>-12600, --- -0.76904296875 + j-0.639099121094
            im_multiplicator=>-10471
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1237),
            data_im_in=>first_stage_im_out(1237),
            product_re_out=>mul_re_out(1237),
            product_im_out=>mul_im_out(1237)
        );

    UMUL_1238 : complex_multiplier
    generic map(
            re_multiplicator=>-13733, --- -0.838195800781 + j-0.545288085938
            im_multiplicator=>-8934
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1238),
            data_im_in=>first_stage_im_out(1238),
            product_re_out=>mul_re_out(1238),
            product_im_out=>mul_im_out(1238)
        );

    UMUL_1239 : complex_multiplier
    generic map(
            re_multiplicator=>-14679, --- -0.895935058594 + j-0.444091796875
            im_multiplicator=>-7276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1239),
            data_im_in=>first_stage_im_out(1239),
            product_re_out=>mul_re_out(1239),
            product_im_out=>mul_im_out(1239)
        );

    UMUL_1240 : complex_multiplier
    generic map(
            re_multiplicator=>-15426, --- -0.941528320312 + j-0.336853027344
            im_multiplicator=>-5519
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1240),
            data_im_in=>first_stage_im_out(1240),
            product_re_out=>mul_re_out(1240),
            product_im_out=>mul_im_out(1240)
        );

    UMUL_1241 : complex_multiplier
    generic map(
            re_multiplicator=>-15963, --- -0.974304199219 + j-0.225036621094
            im_multiplicator=>-3687
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1241),
            data_im_in=>first_stage_im_out(1241),
            product_re_out=>mul_re_out(1241),
            product_im_out=>mul_im_out(1241)
        );

    UMUL_1242 : complex_multiplier
    generic map(
            re_multiplicator=>-16284, --- -0.993896484375 + j-0.110168457031
            im_multiplicator=>-1805
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1242),
            data_im_in=>first_stage_im_out(1242),
            product_re_out=>mul_re_out(1242),
            product_im_out=>mul_im_out(1242)
        );

    UMUL_1243 : complex_multiplier
    generic map(
            re_multiplicator=>-16383, --- -0.999938964844 + j0.006103515625
            im_multiplicator=>100
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1243),
            data_im_in=>first_stage_im_out(1243),
            product_re_out=>mul_re_out(1243),
            product_im_out=>mul_im_out(1243)
        );

    UMUL_1244 : complex_multiplier
    generic map(
            re_multiplicator=>-16260, --- -0.992431640625 + j0.122375488281
            im_multiplicator=>2005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1244),
            data_im_in=>first_stage_im_out(1244),
            product_re_out=>mul_re_out(1244),
            product_im_out=>mul_im_out(1244)
        );

    UMUL_1245 : complex_multiplier
    generic map(
            re_multiplicator=>-15917, --- -0.971496582031 + j0.236999511719
            im_multiplicator=>3883
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1245),
            data_im_in=>first_stage_im_out(1245),
            product_re_out=>mul_re_out(1245),
            product_im_out=>mul_im_out(1245)
        );

    UMUL_1246 : complex_multiplier
    generic map(
            re_multiplicator=>-15357, --- -0.937316894531 + j0.348388671875
            im_multiplicator=>5708
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1246),
            data_im_in=>first_stage_im_out(1246),
            product_re_out=>mul_re_out(1246),
            product_im_out=>mul_im_out(1246)
        );

    UMUL_1247 : complex_multiplier
    generic map(
            re_multiplicator=>-14589, --- -0.890441894531 + j0.455078125
            im_multiplicator=>7456
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1247),
            data_im_in=>first_stage_im_out(1247),
            product_re_out=>mul_re_out(1247),
            product_im_out=>mul_im_out(1247)
        );

    UDELAY_1248_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1248),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1248)
        );
    UDELAY_1248_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1248),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1248)
        );
    USHIFTER_1248_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1248),
            data_out=>mul_re_out(1248)
        );
    USHIFTER_1248_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1248),
            data_out=>mul_im_out(1248)
        );

    UMUL_1249 : complex_multiplier
    generic map(
            re_multiplicator=>16266, --- 0.992797851562 + j-0.119323730469
            im_multiplicator=>-1955
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1249),
            data_im_in=>first_stage_im_out(1249),
            product_re_out=>mul_re_out(1249),
            product_im_out=>mul_im_out(1249)
        );

    UMUL_1250 : complex_multiplier
    generic map(
            re_multiplicator=>15917, --- 0.971496582031 + j-0.236999511719
            im_multiplicator=>-3883
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1250),
            data_im_in=>first_stage_im_out(1250),
            product_re_out=>mul_re_out(1250),
            product_im_out=>mul_im_out(1250)
        );

    UMUL_1251 : complex_multiplier
    generic map(
            re_multiplicator=>15339, --- 0.936218261719 + j-0.351257324219
            im_multiplicator=>-5755
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1251),
            data_im_in=>first_stage_im_out(1251),
            product_re_out=>mul_re_out(1251),
            product_im_out=>mul_im_out(1251)
        );

    UMUL_1252 : complex_multiplier
    generic map(
            re_multiplicator=>14543, --- 0.887634277344 + j-0.460510253906
            im_multiplicator=>-7545
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1252),
            data_im_in=>first_stage_im_out(1252),
            product_re_out=>mul_re_out(1252),
            product_im_out=>mul_im_out(1252)
        );

    UMUL_1253 : complex_multiplier
    generic map(
            re_multiplicator=>13538, --- 0.826293945312 + j-0.563171386719
            im_multiplicator=>-9227
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1253),
            data_im_in=>first_stage_im_out(1253),
            product_re_out=>mul_re_out(1253),
            product_im_out=>mul_im_out(1253)
        );

    UMUL_1254 : complex_multiplier
    generic map(
            re_multiplicator=>12340, --- 0.753173828125 + j-0.657775878906
            im_multiplicator=>-10777
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1254),
            data_im_in=>first_stage_im_out(1254),
            product_re_out=>mul_re_out(1254),
            product_im_out=>mul_im_out(1254)
        );

    UMUL_1255 : complex_multiplier
    generic map(
            re_multiplicator=>10965, --- 0.669250488281 + j-0.742980957031
            im_multiplicator=>-12173
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1255),
            data_im_in=>first_stage_im_out(1255),
            product_re_out=>mul_re_out(1255),
            product_im_out=>mul_im_out(1255)
        );

    UMUL_1256 : complex_multiplier
    generic map(
            re_multiplicator=>9434, --- 0.575805664062 + j-0.817565917969
            im_multiplicator=>-13395
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1256),
            data_im_in=>first_stage_im_out(1256),
            product_re_out=>mul_re_out(1256),
            product_im_out=>mul_im_out(1256)
        );

    UMUL_1257 : complex_multiplier
    generic map(
            re_multiplicator=>7767, --- 0.474060058594 + j-0.880432128906
            im_multiplicator=>-14425
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1257),
            data_im_in=>first_stage_im_out(1257),
            product_re_out=>mul_re_out(1257),
            product_im_out=>mul_im_out(1257)
        );

    UMUL_1258 : complex_multiplier
    generic map(
            re_multiplicator=>5990, --- 0.365600585938 + j-0.930725097656
            im_multiplicator=>-15249
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1258),
            data_im_in=>first_stage_im_out(1258),
            product_re_out=>mul_re_out(1258),
            product_im_out=>mul_im_out(1258)
        );

    UMUL_1259 : complex_multiplier
    generic map(
            re_multiplicator=>4127, --- 0.251892089844 + j-0.967712402344
            im_multiplicator=>-15855
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1259),
            data_im_in=>first_stage_im_out(1259),
            product_re_out=>mul_re_out(1259),
            product_im_out=>mul_im_out(1259)
        );

    UMUL_1260 : complex_multiplier
    generic map(
            re_multiplicator=>2204, --- 0.134521484375 + j-0.990844726562
            im_multiplicator=>-16234
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1260),
            data_im_in=>first_stage_im_out(1260),
            product_re_out=>mul_re_out(1260),
            product_im_out=>mul_im_out(1260)
        );

    UMUL_1261 : complex_multiplier
    generic map(
            re_multiplicator=>251, --- 0.0153198242188 + j-0.999877929688
            im_multiplicator=>-16382
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1261),
            data_im_in=>first_stage_im_out(1261),
            product_re_out=>mul_re_out(1261),
            product_im_out=>mul_im_out(1261)
        );

    UMUL_1262 : complex_multiplier
    generic map(
            re_multiplicator=>-1705, --- -0.104064941406 + j-0.994506835938
            im_multiplicator=>-16294
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1262),
            data_im_in=>first_stage_im_out(1262),
            product_re_out=>mul_re_out(1262),
            product_im_out=>mul_im_out(1262)
        );

    UMUL_1263 : complex_multiplier
    generic map(
            re_multiplicator=>-3638, --- -0.222045898438 + j-0.974975585938
            im_multiplicator=>-15974
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1263),
            data_im_in=>first_stage_im_out(1263),
            product_re_out=>mul_re_out(1263),
            product_im_out=>mul_im_out(1263)
        );

    UMUL_1264 : complex_multiplier
    generic map(
            re_multiplicator=>-5519, --- -0.336853027344 + j-0.941528320312
            im_multiplicator=>-15426
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1264),
            data_im_in=>first_stage_im_out(1264),
            product_re_out=>mul_re_out(1264),
            product_im_out=>mul_im_out(1264)
        );

    UMUL_1265 : complex_multiplier
    generic map(
            re_multiplicator=>-7321, --- -0.446838378906 + j-0.894592285156
            im_multiplicator=>-14657
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1265),
            data_im_in=>first_stage_im_out(1265),
            product_re_out=>mul_re_out(1265),
            product_im_out=>mul_im_out(1265)
        );

    UMUL_1266 : complex_multiplier
    generic map(
            re_multiplicator=>-9018, --- -0.550415039062 + j-0.834838867188
            im_multiplicator=>-13678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1266),
            data_im_in=>first_stage_im_out(1266),
            product_re_out=>mul_re_out(1266),
            product_im_out=>mul_im_out(1266)
        );

    UMUL_1267 : complex_multiplier
    generic map(
            re_multiplicator=>-10586, --- -0.646118164062 + j-0.76318359375
            im_multiplicator=>-12504
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1267),
            data_im_in=>first_stage_im_out(1267),
            product_re_out=>mul_re_out(1267),
            product_im_out=>mul_im_out(1267)
        );

    UMUL_1268 : complex_multiplier
    generic map(
            re_multiplicator=>-12003, --- -0.732604980469 + j-0.680541992188
            im_multiplicator=>-11150
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1268),
            data_im_in=>first_stage_im_out(1268),
            product_re_out=>mul_re_out(1268),
            product_im_out=>mul_im_out(1268)
        );

    UMUL_1269 : complex_multiplier
    generic map(
            re_multiplicator=>-13249, --- -0.808654785156 + j-0.588256835938
            im_multiplicator=>-9638
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1269),
            data_im_in=>first_stage_im_out(1269),
            product_re_out=>mul_re_out(1269),
            product_im_out=>mul_im_out(1269)
        );

    UMUL_1270 : complex_multiplier
    generic map(
            re_multiplicator=>-14304, --- -0.873046875 + j-0.487548828125
            im_multiplicator=>-7988
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1270),
            data_im_in=>first_stage_im_out(1270),
            product_re_out=>mul_re_out(1270),
            product_im_out=>mul_im_out(1270)
        );

    UMUL_1271 : complex_multiplier
    generic map(
            re_multiplicator=>-15156, --- -0.925048828125 + j-0.379821777344
            im_multiplicator=>-6223
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1271),
            data_im_in=>first_stage_im_out(1271),
            product_re_out=>mul_re_out(1271),
            product_im_out=>mul_im_out(1271)
        );

    UMUL_1272 : complex_multiplier
    generic map(
            re_multiplicator=>-15790, --- -0.963745117188 + j-0.266662597656
            im_multiplicator=>-4369
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1272),
            data_im_in=>first_stage_im_out(1272),
            product_re_out=>mul_re_out(1272),
            product_im_out=>mul_im_out(1272)
        );

    UMUL_1273 : complex_multiplier
    generic map(
            re_multiplicator=>-16199, --- -0.988708496094 + j-0.149719238281
            im_multiplicator=>-2453
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1273),
            data_im_in=>first_stage_im_out(1273),
            product_re_out=>mul_re_out(1273),
            product_im_out=>mul_im_out(1273)
        );

    UMUL_1274 : complex_multiplier
    generic map(
            re_multiplicator=>-16376, --- -0.99951171875 + j-0.0306396484375
            im_multiplicator=>-502
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1274),
            data_im_in=>first_stage_im_out(1274),
            product_re_out=>mul_re_out(1274),
            product_im_out=>mul_im_out(1274)
        );

    UMUL_1275 : complex_multiplier
    generic map(
            re_multiplicator=>-16319, --- -0.996032714844 + j0.0888061523438
            im_multiplicator=>1455
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1275),
            data_im_in=>first_stage_im_out(1275),
            product_re_out=>mul_re_out(1275),
            product_im_out=>mul_im_out(1275)
        );

    UMUL_1276 : complex_multiplier
    generic map(
            re_multiplicator=>-16028, --- -0.978271484375 + j0.207092285156
            im_multiplicator=>3393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1276),
            data_im_in=>first_stage_im_out(1276),
            product_re_out=>mul_re_out(1276),
            product_im_out=>mul_im_out(1276)
        );

    UMUL_1277 : complex_multiplier
    generic map(
            re_multiplicator=>-15509, --- -0.946594238281 + j0.322387695312
            im_multiplicator=>5282
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1277),
            data_im_in=>first_stage_im_out(1277),
            product_re_out=>mul_re_out(1277),
            product_im_out=>mul_im_out(1277)
        );

    UMUL_1278 : complex_multiplier
    generic map(
            re_multiplicator=>-14767, --- -0.901306152344 + j0.433044433594
            im_multiplicator=>7095
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1278),
            data_im_in=>first_stage_im_out(1278),
            product_re_out=>mul_re_out(1278),
            product_im_out=>mul_im_out(1278)
        );

    UMUL_1279 : complex_multiplier
    generic map(
            re_multiplicator=>-13815, --- -0.843200683594 + j0.537536621094
            im_multiplicator=>8807
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1279),
            data_im_in=>first_stage_im_out(1279),
            product_re_out=>mul_re_out(1279),
            product_im_out=>mul_im_out(1279)
        );

    UDELAY_1280_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1280),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1280)
        );
    UDELAY_1280_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1280),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1280)
        );
    USHIFTER_1280_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1280),
            data_out=>mul_re_out(1280)
        );
    USHIFTER_1280_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1280),
            data_out=>mul_im_out(1280)
        );

    UMUL_1281 : complex_multiplier
    generic map(
            re_multiplicator=>16260, --- 0.992431640625 + j-0.122375488281
            im_multiplicator=>-2005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1281),
            data_im_in=>first_stage_im_out(1281),
            product_re_out=>mul_re_out(1281),
            product_im_out=>mul_im_out(1281)
        );

    UMUL_1282 : complex_multiplier
    generic map(
            re_multiplicator=>15892, --- 0.969970703125 + j-0.242919921875
            im_multiplicator=>-3980
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1282),
            data_im_in=>first_stage_im_out(1282),
            product_re_out=>mul_re_out(1282),
            product_im_out=>mul_im_out(1282)
        );

    UMUL_1283 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1283),
            data_im_in=>first_stage_im_out(1283),
            product_re_out=>mul_re_out(1283),
            product_im_out=>mul_im_out(1283)
        );

    UMUL_1284 : complex_multiplier
    generic map(
            re_multiplicator=>14449, --- 0.881896972656 + j-0.471374511719
            im_multiplicator=>-7723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1284),
            data_im_in=>first_stage_im_out(1284),
            product_re_out=>mul_re_out(1284),
            product_im_out=>mul_im_out(1284)
        );

    UMUL_1285 : complex_multiplier
    generic map(
            re_multiplicator=>13395, --- 0.817565917969 + j-0.575805664062
            im_multiplicator=>-9434
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1285),
            data_im_in=>first_stage_im_out(1285),
            product_re_out=>mul_re_out(1285),
            product_im_out=>mul_im_out(1285)
        );

    UMUL_1286 : complex_multiplier
    generic map(
            re_multiplicator=>12139, --- 0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1286),
            data_im_in=>first_stage_im_out(1286),
            product_re_out=>mul_re_out(1286),
            product_im_out=>mul_im_out(1286)
        );

    UMUL_1287 : complex_multiplier
    generic map(
            re_multiplicator=>10701, --- 0.653137207031 + j-0.757202148438
            im_multiplicator=>-12406
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1287),
            data_im_in=>first_stage_im_out(1287),
            product_re_out=>mul_re_out(1287),
            product_im_out=>mul_im_out(1287)
        );

    UMUL_1288 : complex_multiplier
    generic map(
            re_multiplicator=>9102, --- 0.555541992188 + j-0.831420898438
            im_multiplicator=>-13622
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1288),
            data_im_in=>first_stage_im_out(1288),
            product_re_out=>mul_re_out(1288),
            product_im_out=>mul_im_out(1288)
        );

    UMUL_1289 : complex_multiplier
    generic map(
            re_multiplicator=>7366, --- 0.449584960938 + j-0.893188476562
            im_multiplicator=>-14634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1289),
            data_im_in=>first_stage_im_out(1289),
            product_re_out=>mul_re_out(1289),
            product_im_out=>mul_im_out(1289)
        );

    UMUL_1290 : complex_multiplier
    generic map(
            re_multiplicator=>5519, --- 0.336853027344 + j-0.941528320312
            im_multiplicator=>-15426
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1290),
            data_im_in=>first_stage_im_out(1290),
            product_re_out=>mul_re_out(1290),
            product_im_out=>mul_im_out(1290)
        );

    UMUL_1291 : complex_multiplier
    generic map(
            re_multiplicator=>3589, --- 0.219055175781 + j-0.975646972656
            im_multiplicator=>-15985
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1291),
            data_im_in=>first_stage_im_out(1291),
            product_re_out=>mul_re_out(1291),
            product_im_out=>mul_im_out(1291)
        );

    UMUL_1292 : complex_multiplier
    generic map(
            re_multiplicator=>1605, --- 0.0979614257812 + j-0.995178222656
            im_multiplicator=>-16305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1292),
            data_im_in=>first_stage_im_out(1292),
            product_re_out=>mul_re_out(1292),
            product_im_out=>mul_im_out(1292)
        );

    UMUL_1293 : complex_multiplier
    generic map(
            re_multiplicator=>-402, --- -0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1293),
            data_im_in=>first_stage_im_out(1293),
            product_re_out=>mul_re_out(1293),
            product_im_out=>mul_im_out(1293)
        );

    UMUL_1294 : complex_multiplier
    generic map(
            re_multiplicator=>-2404, --- -0.146728515625 + j-0.989135742188
            im_multiplicator=>-16206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1294),
            data_im_in=>first_stage_im_out(1294),
            product_re_out=>mul_re_out(1294),
            product_im_out=>mul_im_out(1294)
        );

    UMUL_1295 : complex_multiplier
    generic map(
            re_multiplicator=>-4369, --- -0.266662597656 + j-0.963745117188
            im_multiplicator=>-15790
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1295),
            data_im_in=>first_stage_im_out(1295),
            product_re_out=>mul_re_out(1295),
            product_im_out=>mul_im_out(1295)
        );

    UMUL_1296 : complex_multiplier
    generic map(
            re_multiplicator=>-6269, --- -0.382629394531 + j-0.923828125
            im_multiplicator=>-15136
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1296),
            data_im_in=>first_stage_im_out(1296),
            product_re_out=>mul_re_out(1296),
            product_im_out=>mul_im_out(1296)
        );

    UMUL_1297 : complex_multiplier
    generic map(
            re_multiplicator=>-8075, --- -0.492858886719 + j-0.870056152344
            im_multiplicator=>-14255
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1297),
            data_im_in=>first_stage_im_out(1297),
            product_re_out=>mul_re_out(1297),
            product_im_out=>mul_im_out(1297)
        );

    UMUL_1298 : complex_multiplier
    generic map(
            re_multiplicator=>-9759, --- -0.595642089844 + j-0.803161621094
            im_multiplicator=>-13159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1298),
            data_im_in=>first_stage_im_out(1298),
            product_re_out=>mul_re_out(1298),
            product_im_out=>mul_im_out(1298)
        );

    UMUL_1299 : complex_multiplier
    generic map(
            re_multiplicator=>-11297, --- -0.689514160156 + j-0.724243164062
            im_multiplicator=>-11866
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1299),
            data_im_in=>first_stage_im_out(1299),
            product_re_out=>mul_re_out(1299),
            product_im_out=>mul_im_out(1299)
        );

    UMUL_1300 : complex_multiplier
    generic map(
            re_multiplicator=>-12665, --- -0.773010253906 + j-0.634338378906
            im_multiplicator=>-10393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1300),
            data_im_in=>first_stage_im_out(1300),
            product_re_out=>mul_re_out(1300),
            product_im_out=>mul_im_out(1300)
        );

    UMUL_1301 : complex_multiplier
    generic map(
            re_multiplicator=>-13842, --- -0.844848632812 + j-0.534973144531
            im_multiplicator=>-8765
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1301),
            data_im_in=>first_stage_im_out(1301),
            product_re_out=>mul_re_out(1301),
            product_im_out=>mul_im_out(1301)
        );

    UMUL_1302 : complex_multiplier
    generic map(
            re_multiplicator=>-14810, --- -0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1302),
            data_im_in=>first_stage_im_out(1302),
            product_re_out=>mul_re_out(1302),
            product_im_out=>mul_im_out(1302)
        );

    UMUL_1303 : complex_multiplier
    generic map(
            re_multiplicator=>-15557, --- -0.949523925781 + j-0.313659667969
            im_multiplicator=>-5139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1303),
            data_im_in=>first_stage_im_out(1303),
            product_re_out=>mul_re_out(1303),
            product_im_out=>mul_im_out(1303)
        );

    UMUL_1304 : complex_multiplier
    generic map(
            re_multiplicator=>-16069, --- -0.980773925781 + j-0.195068359375
            im_multiplicator=>-3196
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1304),
            data_im_in=>first_stage_im_out(1304),
            product_re_out=>mul_re_out(1304),
            product_im_out=>mul_im_out(1304)
        );

    UMUL_1305 : complex_multiplier
    generic map(
            re_multiplicator=>-16339, --- -0.997253417969 + j-0.0735473632812
            im_multiplicator=>-1205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1305),
            data_im_in=>first_stage_im_out(1305),
            product_re_out=>mul_re_out(1305),
            product_im_out=>mul_im_out(1305)
        );

    UMUL_1306 : complex_multiplier
    generic map(
            re_multiplicator=>-16364, --- -0.998779296875 + j0.0490112304688
            im_multiplicator=>803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1306),
            data_im_in=>first_stage_im_out(1306),
            product_re_out=>mul_re_out(1306),
            product_im_out=>mul_im_out(1306)
        );

    UMUL_1307 : complex_multiplier
    generic map(
            re_multiplicator=>-16142, --- -0.985229492188 + j0.170959472656
            im_multiplicator=>2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1307),
            data_im_in=>first_stage_im_out(1307),
            product_re_out=>mul_re_out(1307),
            product_im_out=>mul_im_out(1307)
        );

    UMUL_1308 : complex_multiplier
    generic map(
            re_multiplicator=>-15678, --- -0.956909179688 + j0.290283203125
            im_multiplicator=>4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1308),
            data_im_in=>first_stage_im_out(1308),
            product_re_out=>mul_re_out(1308),
            product_im_out=>mul_im_out(1308)
        );

    UMUL_1309 : complex_multiplier
    generic map(
            re_multiplicator=>-14978, --- -0.914184570312 + j0.405212402344
            im_multiplicator=>6639
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1309),
            data_im_in=>first_stage_im_out(1309),
            product_re_out=>mul_re_out(1309),
            product_im_out=>mul_im_out(1309)
        );

    UMUL_1310 : complex_multiplier
    generic map(
            re_multiplicator=>-14053, --- -0.857727050781 + j0.514099121094
            im_multiplicator=>8423
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1310),
            data_im_in=>first_stage_im_out(1310),
            product_re_out=>mul_re_out(1310),
            product_im_out=>mul_im_out(1310)
        );

    UMUL_1311 : complex_multiplier
    generic map(
            re_multiplicator=>-12916, --- -0.788330078125 + j0.615173339844
            im_multiplicator=>10079
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1311),
            data_im_in=>first_stage_im_out(1311),
            product_re_out=>mul_re_out(1311),
            product_im_out=>mul_im_out(1311)
        );

    UDELAY_1312_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1312),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1312)
        );
    UDELAY_1312_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1312),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1312)
        );
    USHIFTER_1312_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1312),
            data_out=>mul_re_out(1312)
        );
    USHIFTER_1312_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1312),
            data_out=>mul_im_out(1312)
        );

    UMUL_1313 : complex_multiplier
    generic map(
            re_multiplicator=>16254, --- 0.992065429688 + j-0.125427246094
            im_multiplicator=>-2055
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1313),
            data_im_in=>first_stage_im_out(1313),
            product_re_out=>mul_re_out(1313),
            product_im_out=>mul_im_out(1313)
        );

    UMUL_1314 : complex_multiplier
    generic map(
            re_multiplicator=>15868, --- 0.968505859375 + j-0.248901367188
            im_multiplicator=>-4078
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1314),
            data_im_in=>first_stage_im_out(1314),
            product_re_out=>mul_re_out(1314),
            product_im_out=>mul_im_out(1314)
        );

    UMUL_1315 : complex_multiplier
    generic map(
            re_multiplicator=>15231, --- 0.929626464844 + j-0.368408203125
            im_multiplicator=>-6036
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1315),
            data_im_in=>first_stage_im_out(1315),
            product_re_out=>mul_re_out(1315),
            product_im_out=>mul_im_out(1315)
        );

    UMUL_1316 : complex_multiplier
    generic map(
            re_multiplicator=>14353, --- 0.876037597656 + j-0.482177734375
            im_multiplicator=>-7900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1316),
            data_im_in=>first_stage_im_out(1316),
            product_re_out=>mul_re_out(1316),
            product_im_out=>mul_im_out(1316)
        );

    UMUL_1317 : complex_multiplier
    generic map(
            re_multiplicator=>13249, --- 0.808654785156 + j-0.588256835938
            im_multiplicator=>-9638
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1317),
            data_im_in=>first_stage_im_out(1317),
            product_re_out=>mul_re_out(1317),
            product_im_out=>mul_im_out(1317)
        );

    UMUL_1318 : complex_multiplier
    generic map(
            re_multiplicator=>11935, --- 0.728454589844 + j-0.68505859375
            im_multiplicator=>-11224
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1318),
            data_im_in=>first_stage_im_out(1318),
            product_re_out=>mul_re_out(1318),
            product_im_out=>mul_im_out(1318)
        );

    UMUL_1319 : complex_multiplier
    generic map(
            re_multiplicator=>10432, --- 0.63671875 + j-0.771057128906
            im_multiplicator=>-12633
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1319),
            data_im_in=>first_stage_im_out(1319),
            product_re_out=>mul_re_out(1319),
            product_im_out=>mul_im_out(1319)
        );

    UMUL_1320 : complex_multiplier
    generic map(
            re_multiplicator=>8765, --- 0.534973144531 + j-0.844848632812
            im_multiplicator=>-13842
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1320),
            data_im_in=>first_stage_im_out(1320),
            product_re_out=>mul_re_out(1320),
            product_im_out=>mul_im_out(1320)
        );

    UMUL_1321 : complex_multiplier
    generic map(
            re_multiplicator=>6959, --- 0.424743652344 + j-0.9052734375
            im_multiplicator=>-14832
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1321),
            data_im_in=>first_stage_im_out(1321),
            product_re_out=>mul_re_out(1321),
            product_im_out=>mul_im_out(1321)
        );

    UMUL_1322 : complex_multiplier
    generic map(
            re_multiplicator=>5043, --- 0.307800292969 + j-0.951416015625
            im_multiplicator=>-15588
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1322),
            data_im_in=>first_stage_im_out(1322),
            product_re_out=>mul_re_out(1322),
            product_im_out=>mul_im_out(1322)
        );

    UMUL_1323 : complex_multiplier
    generic map(
            re_multiplicator=>3048, --- 0.18603515625 + j-0.982482910156
            im_multiplicator=>-16097
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1323),
            data_im_in=>first_stage_im_out(1323),
            product_re_out=>mul_re_out(1323),
            product_im_out=>mul_im_out(1323)
        );

    UMUL_1324 : complex_multiplier
    generic map(
            re_multiplicator=>1004, --- 0.061279296875 + j-0.998107910156
            im_multiplicator=>-16353
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1324),
            data_im_in=>first_stage_im_out(1324),
            product_re_out=>mul_re_out(1324),
            product_im_out=>mul_im_out(1324)
        );

    UMUL_1325 : complex_multiplier
    generic map(
            re_multiplicator=>-1054, --- -0.0643310546875 + j-0.997924804688
            im_multiplicator=>-16350
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1325),
            data_im_in=>first_stage_im_out(1325),
            product_re_out=>mul_re_out(1325),
            product_im_out=>mul_im_out(1325)
        );

    UMUL_1326 : complex_multiplier
    generic map(
            re_multiplicator=>-3097, --- -0.189025878906 + j-0.98193359375
            im_multiplicator=>-16088
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1326),
            data_im_in=>first_stage_im_out(1326),
            product_re_out=>mul_re_out(1326),
            product_im_out=>mul_im_out(1326)
        );

    UMUL_1327 : complex_multiplier
    generic map(
            re_multiplicator=>-5091, --- -0.310729980469 + j-0.950439453125
            im_multiplicator=>-15572
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1327),
            data_im_in=>first_stage_im_out(1327),
            product_re_out=>mul_re_out(1327),
            product_im_out=>mul_im_out(1327)
        );

    UMUL_1328 : complex_multiplier
    generic map(
            re_multiplicator=>-7005, --- -0.427551269531 + j-0.903930664062
            im_multiplicator=>-14810
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1328),
            data_im_in=>first_stage_im_out(1328),
            product_re_out=>mul_re_out(1328),
            product_im_out=>mul_im_out(1328)
        );

    UMUL_1329 : complex_multiplier
    generic map(
            re_multiplicator=>-8807, --- -0.537536621094 + j-0.843200683594
            im_multiplicator=>-13815
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1329),
            data_im_in=>first_stage_im_out(1329),
            product_re_out=>mul_re_out(1329),
            product_im_out=>mul_im_out(1329)
        );

    UMUL_1330 : complex_multiplier
    generic map(
            re_multiplicator=>-10471, --- -0.639099121094 + j-0.76904296875
            im_multiplicator=>-12600
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1330),
            data_im_in=>first_stage_im_out(1330),
            product_re_out=>mul_re_out(1330),
            product_im_out=>mul_im_out(1330)
        );

    UMUL_1331 : complex_multiplier
    generic map(
            re_multiplicator=>-11969, --- -0.730529785156 + j-0.682800292969
            im_multiplicator=>-11187
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1331),
            data_im_in=>first_stage_im_out(1331),
            product_re_out=>mul_re_out(1331),
            product_im_out=>mul_im_out(1331)
        );

    UMUL_1332 : complex_multiplier
    generic map(
            re_multiplicator=>-13278, --- -0.810424804688 + j-0.585754394531
            im_multiplicator=>-9597
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1332),
            data_im_in=>first_stage_im_out(1332),
            product_re_out=>mul_re_out(1332),
            product_im_out=>mul_im_out(1332)
        );

    UMUL_1333 : complex_multiplier
    generic map(
            re_multiplicator=>-14377, --- -0.877502441406 + j-0.4794921875
            im_multiplicator=>-7856
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1333),
            data_im_in=>first_stage_im_out(1333),
            product_re_out=>mul_re_out(1333),
            product_im_out=>mul_im_out(1333)
        );

    UMUL_1334 : complex_multiplier
    generic map(
            re_multiplicator=>-15249, --- -0.930725097656 + j-0.365600585938
            im_multiplicator=>-5990
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1334),
            data_im_in=>first_stage_im_out(1334),
            product_re_out=>mul_re_out(1334),
            product_im_out=>mul_im_out(1334)
        );

    UMUL_1335 : complex_multiplier
    generic map(
            re_multiplicator=>-15880, --- -0.96923828125 + j-0.245910644531
            im_multiplicator=>-4029
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1335),
            data_im_in=>first_stage_im_out(1335),
            product_re_out=>mul_re_out(1335),
            product_im_out=>mul_im_out(1335)
        );

    UMUL_1336 : complex_multiplier
    generic map(
            re_multiplicator=>-16260, --- -0.992431640625 + j-0.122375488281
            im_multiplicator=>-2005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1336),
            data_im_in=>first_stage_im_out(1336),
            product_re_out=>mul_re_out(1336),
            product_im_out=>mul_im_out(1336)
        );

    UMUL_1337 : complex_multiplier
    generic map(
            re_multiplicator=>-16383, --- -0.999938964844 + j0.0030517578125
            im_multiplicator=>50
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1337),
            data_im_in=>first_stage_im_out(1337),
            product_re_out=>mul_re_out(1337),
            product_im_out=>mul_im_out(1337)
        );

    UMUL_1338 : complex_multiplier
    generic map(
            re_multiplicator=>-16248, --- -0.99169921875 + j0.128479003906
            im_multiplicator=>2105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1338),
            data_im_in=>first_stage_im_out(1338),
            product_re_out=>mul_re_out(1338),
            product_im_out=>mul_im_out(1338)
        );

    UMUL_1339 : complex_multiplier
    generic map(
            re_multiplicator=>-15855, --- -0.967712402344 + j0.251892089844
            im_multiplicator=>4127
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1339),
            data_im_in=>first_stage_im_out(1339),
            product_re_out=>mul_re_out(1339),
            product_im_out=>mul_im_out(1339)
        );

    UMUL_1340 : complex_multiplier
    generic map(
            re_multiplicator=>-15212, --- -0.928466796875 + j0.371276855469
            im_multiplicator=>6083
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1340),
            data_im_in=>first_stage_im_out(1340),
            product_re_out=>mul_re_out(1340),
            product_im_out=>mul_im_out(1340)
        );

    UMUL_1341 : complex_multiplier
    generic map(
            re_multiplicator=>-14329, --- -0.874572753906 + j0.48486328125
            im_multiplicator=>7944
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1341),
            data_im_in=>first_stage_im_out(1341),
            product_re_out=>mul_re_out(1341),
            product_im_out=>mul_im_out(1341)
        );

    UMUL_1342 : complex_multiplier
    generic map(
            re_multiplicator=>-13219, --- -0.806823730469 + j0.590759277344
            im_multiplicator=>9679
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1342),
            data_im_in=>first_stage_im_out(1342),
            product_re_out=>mul_re_out(1342),
            product_im_out=>mul_im_out(1342)
        );

    UMUL_1343 : complex_multiplier
    generic map(
            re_multiplicator=>-11900, --- -0.726318359375 + j0.687255859375
            im_multiplicator=>11260
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1343),
            data_im_in=>first_stage_im_out(1343),
            product_re_out=>mul_re_out(1343),
            product_im_out=>mul_im_out(1343)
        );

    UDELAY_1344_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1344),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1344)
        );
    UDELAY_1344_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1344),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1344)
        );
    USHIFTER_1344_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1344),
            data_out=>mul_re_out(1344)
        );
    USHIFTER_1344_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1344),
            data_out=>mul_im_out(1344)
        );

    UMUL_1345 : complex_multiplier
    generic map(
            re_multiplicator=>16248, --- 0.99169921875 + j-0.128479003906
            im_multiplicator=>-2105
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1345),
            data_im_in=>first_stage_im_out(1345),
            product_re_out=>mul_re_out(1345),
            product_im_out=>mul_im_out(1345)
        );

    UMUL_1346 : complex_multiplier
    generic map(
            re_multiplicator=>15842, --- 0.966918945312 + j-0.254821777344
            im_multiplicator=>-4175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1346),
            data_im_in=>first_stage_im_out(1346),
            product_re_out=>mul_re_out(1346),
            product_im_out=>mul_im_out(1346)
        );

    UMUL_1347 : complex_multiplier
    generic map(
            re_multiplicator=>15175, --- 0.926208496094 + j-0.376953125
            im_multiplicator=>-6176
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1347),
            data_im_in=>first_stage_im_out(1347),
            product_re_out=>mul_re_out(1347),
            product_im_out=>mul_im_out(1347)
        );

    UMUL_1348 : complex_multiplier
    generic map(
            re_multiplicator=>14255, --- 0.870056152344 + j-0.492858886719
            im_multiplicator=>-8075
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1348),
            data_im_in=>first_stage_im_out(1348),
            product_re_out=>mul_re_out(1348),
            product_im_out=>mul_im_out(1348)
        );

    UMUL_1349 : complex_multiplier
    generic map(
            re_multiplicator=>13099, --- 0.799499511719 + j-0.6005859375
            im_multiplicator=>-9840
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1349),
            data_im_in=>first_stage_im_out(1349),
            product_re_out=>mul_re_out(1349),
            product_im_out=>mul_im_out(1349)
        );

    UMUL_1350 : complex_multiplier
    generic map(
            re_multiplicator=>11726, --- 0.715698242188 + j-0.698364257812
            im_multiplicator=>-11442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1350),
            data_im_in=>first_stage_im_out(1350),
            product_re_out=>mul_re_out(1350),
            product_im_out=>mul_im_out(1350)
        );

    UMUL_1351 : complex_multiplier
    generic map(
            re_multiplicator=>10159, --- 0.620056152344 + j-0.784545898438
            im_multiplicator=>-12854
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1351),
            data_im_in=>first_stage_im_out(1351),
            product_re_out=>mul_re_out(1351),
            product_im_out=>mul_im_out(1351)
        );

    UMUL_1352 : complex_multiplier
    generic map(
            re_multiplicator=>8423, --- 0.514099121094 + j-0.857727050781
            im_multiplicator=>-14053
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1352),
            data_im_in=>first_stage_im_out(1352),
            product_re_out=>mul_re_out(1352),
            product_im_out=>mul_im_out(1352)
        );

    UMUL_1353 : complex_multiplier
    generic map(
            re_multiplicator=>6547, --- 0.399597167969 + j-0.916625976562
            im_multiplicator=>-15018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1353),
            data_im_in=>first_stage_im_out(1353),
            product_re_out=>mul_re_out(1353),
            product_im_out=>mul_im_out(1353)
        );

    UMUL_1354 : complex_multiplier
    generic map(
            re_multiplicator=>4563, --- 0.278503417969 + j-0.960388183594
            im_multiplicator=>-15735
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1354),
            data_im_in=>first_stage_im_out(1354),
            product_re_out=>mul_re_out(1354),
            product_im_out=>mul_im_out(1354)
        );

    UMUL_1355 : complex_multiplier
    generic map(
            re_multiplicator=>2503, --- 0.152770996094 + j-0.988220214844
            im_multiplicator=>-16191
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1355),
            data_im_in=>first_stage_im_out(1355),
            product_re_out=>mul_re_out(1355),
            product_im_out=>mul_im_out(1355)
        );

    UMUL_1356 : complex_multiplier
    generic map(
            re_multiplicator=>402, --- 0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1356),
            data_im_in=>first_stage_im_out(1356),
            product_re_out=>mul_re_out(1356),
            product_im_out=>mul_im_out(1356)
        );

    UMUL_1357 : complex_multiplier
    generic map(
            re_multiplicator=>-1705, --- -0.104064941406 + j-0.994506835938
            im_multiplicator=>-16294
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1357),
            data_im_in=>first_stage_im_out(1357),
            product_re_out=>mul_re_out(1357),
            product_im_out=>mul_im_out(1357)
        );

    UMUL_1358 : complex_multiplier
    generic map(
            re_multiplicator=>-3785, --- -0.231018066406 + j-0.972900390625
            im_multiplicator=>-15940
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1358),
            data_im_in=>first_stage_im_out(1358),
            product_re_out=>mul_re_out(1358),
            product_im_out=>mul_im_out(1358)
        );

    UMUL_1359 : complex_multiplier
    generic map(
            re_multiplicator=>-5802, --- -0.354125976562 + j-0.935180664062
            im_multiplicator=>-15322
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1359),
            data_im_in=>first_stage_im_out(1359),
            product_re_out=>mul_re_out(1359),
            product_im_out=>mul_im_out(1359)
        );

    UMUL_1360 : complex_multiplier
    generic map(
            re_multiplicator=>-7723, --- -0.471374511719 + j-0.881896972656
            im_multiplicator=>-14449
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1360),
            data_im_in=>first_stage_im_out(1360),
            product_re_out=>mul_re_out(1360),
            product_im_out=>mul_im_out(1360)
        );

    UMUL_1361 : complex_multiplier
    generic map(
            re_multiplicator=>-9516, --- -0.580810546875 + j-0.814025878906
            im_multiplicator=>-13337
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1361),
            data_im_in=>first_stage_im_out(1361),
            product_re_out=>mul_re_out(1361),
            product_im_out=>mul_im_out(1361)
        );

    UMUL_1362 : complex_multiplier
    generic map(
            re_multiplicator=>-11150, --- -0.680541992188 + j-0.732604980469
            im_multiplicator=>-12003
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1362),
            data_im_in=>first_stage_im_out(1362),
            product_re_out=>mul_re_out(1362),
            product_im_out=>mul_im_out(1362)
        );

    UMUL_1363 : complex_multiplier
    generic map(
            re_multiplicator=>-12600, --- -0.76904296875 + j-0.639099121094
            im_multiplicator=>-10471
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1363),
            data_im_in=>first_stage_im_out(1363),
            product_re_out=>mul_re_out(1363),
            product_im_out=>mul_im_out(1363)
        );

    UMUL_1364 : complex_multiplier
    generic map(
            re_multiplicator=>-13842, --- -0.844848632812 + j-0.534973144531
            im_multiplicator=>-8765
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1364),
            data_im_in=>first_stage_im_out(1364),
            product_re_out=>mul_re_out(1364),
            product_im_out=>mul_im_out(1364)
        );

    UMUL_1365 : complex_multiplier
    generic map(
            re_multiplicator=>-14853, --- -0.906555175781 + j-0.421997070312
            im_multiplicator=>-6914
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1365),
            data_im_in=>first_stage_im_out(1365),
            product_re_out=>mul_re_out(1365),
            product_im_out=>mul_im_out(1365)
        );

    UMUL_1366 : complex_multiplier
    generic map(
            re_multiplicator=>-15618, --- -0.953247070312 + j-0.302001953125
            im_multiplicator=>-4948
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1366),
            data_im_in=>first_stage_im_out(1366),
            product_re_out=>mul_re_out(1366),
            product_im_out=>mul_im_out(1366)
        );

    UMUL_1367 : complex_multiplier
    generic map(
            re_multiplicator=>-16125, --- -0.984191894531 + j-0.177001953125
            im_multiplicator=>-2900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1367),
            data_im_in=>first_stage_im_out(1367),
            product_re_out=>mul_re_out(1367),
            product_im_out=>mul_im_out(1367)
        );

    UMUL_1368 : complex_multiplier
    generic map(
            re_multiplicator=>-16364, --- -0.998779296875 + j-0.0490112304688
            im_multiplicator=>-803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1368),
            data_im_in=>first_stage_im_out(1368),
            product_re_out=>mul_re_out(1368),
            product_im_out=>mul_im_out(1368)
        );

    UMUL_1369 : complex_multiplier
    generic map(
            re_multiplicator=>-16331, --- -0.996765136719 + j0.0796508789062
            im_multiplicator=>1305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1369),
            data_im_in=>first_stage_im_out(1369),
            product_re_out=>mul_re_out(1369),
            product_im_out=>mul_im_out(1369)
        );

    UMUL_1370 : complex_multiplier
    generic map(
            re_multiplicator=>-16028, --- -0.978271484375 + j0.207092285156
            im_multiplicator=>3393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1370),
            data_im_in=>first_stage_im_out(1370),
            product_re_out=>mul_re_out(1370),
            product_im_out=>mul_im_out(1370)
        );

    UMUL_1371 : complex_multiplier
    generic map(
            re_multiplicator=>-15459, --- -0.943542480469 + j0.3310546875
            im_multiplicator=>5424
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1371),
            data_im_in=>first_stage_im_out(1371),
            product_re_out=>mul_re_out(1371),
            product_im_out=>mul_im_out(1371)
        );

    UMUL_1372 : complex_multiplier
    generic map(
            re_multiplicator=>-14634, --- -0.893188476562 + j0.449584960938
            im_multiplicator=>7366
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1372),
            data_im_in=>first_stage_im_out(1372),
            product_re_out=>mul_re_out(1372),
            product_im_out=>mul_im_out(1372)
        );

    UMUL_1373 : complex_multiplier
    generic map(
            re_multiplicator=>-13566, --- -0.828002929688 + j0.560607910156
            im_multiplicator=>9185
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1373),
            data_im_in=>first_stage_im_out(1373),
            product_re_out=>mul_re_out(1373),
            product_im_out=>mul_im_out(1373)
        );

    UMUL_1374 : complex_multiplier
    generic map(
            re_multiplicator=>-12273, --- -0.749084472656 + j0.662414550781
            im_multiplicator=>10853
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1374),
            data_im_in=>first_stage_im_out(1374),
            product_re_out=>mul_re_out(1374),
            product_im_out=>mul_im_out(1374)
        );

    UMUL_1375 : complex_multiplier
    generic map(
            re_multiplicator=>-10777, --- -0.657775878906 + j0.753173828125
            im_multiplicator=>12340
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1375),
            data_im_in=>first_stage_im_out(1375),
            product_re_out=>mul_re_out(1375),
            product_im_out=>mul_im_out(1375)
        );

    UDELAY_1376_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1376),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1376)
        );
    UDELAY_1376_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1376),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1376)
        );
    USHIFTER_1376_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1376),
            data_out=>mul_re_out(1376)
        );
    USHIFTER_1376_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1376),
            data_out=>mul_im_out(1376)
        );

    UMUL_1377 : complex_multiplier
    generic map(
            re_multiplicator=>16241, --- 0.991271972656 + j-0.131530761719
            im_multiplicator=>-2155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1377),
            data_im_in=>first_stage_im_out(1377),
            product_re_out=>mul_re_out(1377),
            product_im_out=>mul_im_out(1377)
        );

    UMUL_1378 : complex_multiplier
    generic map(
            re_multiplicator=>15817, --- 0.965393066406 + j-0.2607421875
            im_multiplicator=>-4272
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1378),
            data_im_in=>first_stage_im_out(1378),
            product_re_out=>mul_re_out(1378),
            product_im_out=>mul_im_out(1378)
        );

    UMUL_1379 : complex_multiplier
    generic map(
            re_multiplicator=>15117, --- 0.922668457031 + j-0.385498046875
            im_multiplicator=>-6316
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1379),
            data_im_in=>first_stage_im_out(1379),
            product_re_out=>mul_re_out(1379),
            product_im_out=>mul_im_out(1379)
        );

    UMUL_1380 : complex_multiplier
    generic map(
            re_multiplicator=>14155, --- 0.863952636719 + j-0.503479003906
            im_multiplicator=>-8249
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1380),
            data_im_in=>first_stage_im_out(1380),
            product_re_out=>mul_re_out(1380),
            product_im_out=>mul_im_out(1380)
        );

    UMUL_1381 : complex_multiplier
    generic map(
            re_multiplicator=>12947, --- 0.790222167969 + j-0.61279296875
            im_multiplicator=>-10040
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1381),
            data_im_in=>first_stage_im_out(1381),
            product_re_out=>mul_re_out(1381),
            product_im_out=>mul_im_out(1381)
        );

    UMUL_1382 : complex_multiplier
    generic map(
            re_multiplicator=>11513, --- 0.702697753906 + j-0.71142578125
            im_multiplicator=>-11656
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1382),
            data_im_in=>first_stage_im_out(1382),
            product_re_out=>mul_re_out(1382),
            product_im_out=>mul_im_out(1382)
        );

    UMUL_1383 : complex_multiplier
    generic map(
            re_multiplicator=>9880, --- 0.60302734375 + j-0.797668457031
            im_multiplicator=>-13069
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1383),
            data_im_in=>first_stage_im_out(1383),
            product_re_out=>mul_re_out(1383),
            product_im_out=>mul_im_out(1383)
        );

    UMUL_1384 : complex_multiplier
    generic map(
            re_multiplicator=>8075, --- 0.492858886719 + j-0.870056152344
            im_multiplicator=>-14255
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1384),
            data_im_in=>first_stage_im_out(1384),
            product_re_out=>mul_re_out(1384),
            product_im_out=>mul_im_out(1384)
        );

    UMUL_1385 : complex_multiplier
    generic map(
            re_multiplicator=>6130, --- 0.374145507812 + j-0.927307128906
            im_multiplicator=>-15193
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1385),
            data_im_in=>first_stage_im_out(1385),
            product_re_out=>mul_re_out(1385),
            product_im_out=>mul_im_out(1385)
        );

    UMUL_1386 : complex_multiplier
    generic map(
            re_multiplicator=>4078, --- 0.248901367188 + j-0.968505859375
            im_multiplicator=>-15868
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1386),
            data_im_in=>first_stage_im_out(1386),
            product_re_out=>mul_re_out(1386),
            product_im_out=>mul_im_out(1386)
        );

    UMUL_1387 : complex_multiplier
    generic map(
            re_multiplicator=>1955, --- 0.119323730469 + j-0.992797851562
            im_multiplicator=>-16266
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1387),
            data_im_in=>first_stage_im_out(1387),
            product_re_out=>mul_re_out(1387),
            product_im_out=>mul_im_out(1387)
        );

    UMUL_1388 : complex_multiplier
    generic map(
            re_multiplicator=>-201, --- -0.0122680664062 + j-0.999877929688
            im_multiplicator=>-16382
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1388),
            data_im_in=>first_stage_im_out(1388),
            product_re_out=>mul_re_out(1388),
            product_im_out=>mul_im_out(1388)
        );

    UMUL_1389 : complex_multiplier
    generic map(
            re_multiplicator=>-2354, --- -0.143676757812 + j-0.989562988281
            im_multiplicator=>-16213
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1389),
            data_im_in=>first_stage_im_out(1389),
            product_re_out=>mul_re_out(1389),
            product_im_out=>mul_im_out(1389)
        );

    UMUL_1390 : complex_multiplier
    generic map(
            re_multiplicator=>-4466, --- -0.272583007812 + j-0.962097167969
            im_multiplicator=>-15763
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1390),
            data_im_in=>first_stage_im_out(1390),
            product_re_out=>mul_re_out(1390),
            product_im_out=>mul_im_out(1390)
        );

    UMUL_1391 : complex_multiplier
    generic map(
            re_multiplicator=>-6501, --- -0.396789550781 + j-0.917846679688
            im_multiplicator=>-15038
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1391),
            data_im_in=>first_stage_im_out(1391),
            product_re_out=>mul_re_out(1391),
            product_im_out=>mul_im_out(1391)
        );

    UMUL_1392 : complex_multiplier
    generic map(
            re_multiplicator=>-8423, --- -0.514099121094 + j-0.857727050781
            im_multiplicator=>-14053
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1392),
            data_im_in=>first_stage_im_out(1392),
            product_re_out=>mul_re_out(1392),
            product_im_out=>mul_im_out(1392)
        );

    UMUL_1393 : complex_multiplier
    generic map(
            re_multiplicator=>-10198, --- -0.622436523438 + j-0.782592773438
            im_multiplicator=>-12822
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1393),
            data_im_in=>first_stage_im_out(1393),
            product_re_out=>mul_re_out(1393),
            product_im_out=>mul_im_out(1393)
        );

    UMUL_1394 : complex_multiplier
    generic map(
            re_multiplicator=>-11796, --- -0.719970703125 + j-0.693969726562
            im_multiplicator=>-11370
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1394),
            data_im_in=>first_stage_im_out(1394),
            product_re_out=>mul_re_out(1394),
            product_im_out=>mul_im_out(1394)
        );

    UMUL_1395 : complex_multiplier
    generic map(
            re_multiplicator=>-13189, --- -0.804992675781 + j-0.593200683594
            im_multiplicator=>-9719
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1395),
            data_im_in=>first_stage_im_out(1395),
            product_re_out=>mul_re_out(1395),
            product_im_out=>mul_im_out(1395)
        );

    UMUL_1396 : complex_multiplier
    generic map(
            re_multiplicator=>-14353, --- -0.876037597656 + j-0.482177734375
            im_multiplicator=>-7900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1396),
            data_im_in=>first_stage_im_out(1396),
            product_re_out=>mul_re_out(1396),
            product_im_out=>mul_im_out(1396)
        );

    UMUL_1397 : complex_multiplier
    generic map(
            re_multiplicator=>-15267, --- -0.931823730469 + j-0.362731933594
            im_multiplicator=>-5943
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1397),
            data_im_in=>first_stage_im_out(1397),
            product_re_out=>mul_re_out(1397),
            product_im_out=>mul_im_out(1397)
        );

    UMUL_1398 : complex_multiplier
    generic map(
            re_multiplicator=>-15917, --- -0.971496582031 + j-0.236999511719
            im_multiplicator=>-3883
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1398),
            data_im_in=>first_stage_im_out(1398),
            product_re_out=>mul_re_out(1398),
            product_im_out=>mul_im_out(1398)
        );

    UMUL_1399 : complex_multiplier
    generic map(
            re_multiplicator=>-16289, --- -0.994201660156 + j-0.107116699219
            im_multiplicator=>-1755
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1399),
            data_im_in=>first_stage_im_out(1399),
            product_re_out=>mul_re_out(1399),
            product_im_out=>mul_im_out(1399)
        );

    UMUL_1400 : complex_multiplier
    generic map(
            re_multiplicator=>-16379, --- -0.999694824219 + j0.0245361328125
            im_multiplicator=>402
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1400),
            data_im_in=>first_stage_im_out(1400),
            product_re_out=>mul_re_out(1400),
            product_im_out=>mul_im_out(1400)
        );

    UMUL_1401 : complex_multiplier
    generic map(
            re_multiplicator=>-16183, --- -0.987731933594 + j0.155822753906
            im_multiplicator=>2553
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1401),
            data_im_in=>first_stage_im_out(1401),
            product_re_out=>mul_re_out(1401),
            product_im_out=>mul_im_out(1401)
        );

    UMUL_1402 : complex_multiplier
    generic map(
            re_multiplicator=>-15707, --- -0.958679199219 + j0.284362792969
            im_multiplicator=>4659
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1402),
            data_im_in=>first_stage_im_out(1402),
            product_re_out=>mul_re_out(1402),
            product_im_out=>mul_im_out(1402)
        );

    UMUL_1403 : complex_multiplier
    generic map(
            re_multiplicator=>-14957, --- -0.912902832031 + j0.408020019531
            im_multiplicator=>6685
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1403),
            data_im_in=>first_stage_im_out(1403),
            product_re_out=>mul_re_out(1403),
            product_im_out=>mul_im_out(1403)
        );

    UMUL_1404 : complex_multiplier
    generic map(
            re_multiplicator=>-13948, --- -0.851318359375 + j0.524536132812
            im_multiplicator=>8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1404),
            data_im_in=>first_stage_im_out(1404),
            product_re_out=>mul_re_out(1404),
            product_im_out=>mul_im_out(1404)
        );

    UMUL_1405 : complex_multiplier
    generic map(
            re_multiplicator=>-12696, --- -0.77490234375 + j0.631958007812
            im_multiplicator=>10354
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1405),
            data_im_in=>first_stage_im_out(1405),
            product_re_out=>mul_re_out(1405),
            product_im_out=>mul_im_out(1405)
        );

    UMUL_1406 : complex_multiplier
    generic map(
            re_multiplicator=>-11224, --- -0.68505859375 + j0.728454589844
            im_multiplicator=>11935
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1406),
            data_im_in=>first_stage_im_out(1406),
            product_re_out=>mul_re_out(1406),
            product_im_out=>mul_im_out(1406)
        );

    UMUL_1407 : complex_multiplier
    generic map(
            re_multiplicator=>-9556, --- -0.583251953125 + j0.812194824219
            im_multiplicator=>13307
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1407),
            data_im_in=>first_stage_im_out(1407),
            product_re_out=>mul_re_out(1407),
            product_im_out=>mul_im_out(1407)
        );

    UDELAY_1408_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1408),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1408)
        );
    UDELAY_1408_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1408),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1408)
        );
    USHIFTER_1408_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1408),
            data_out=>mul_re_out(1408)
        );
    USHIFTER_1408_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1408),
            data_out=>mul_im_out(1408)
        );

    UMUL_1409 : complex_multiplier
    generic map(
            re_multiplicator=>16234, --- 0.990844726562 + j-0.134521484375
            im_multiplicator=>-2204
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1409),
            data_im_in=>first_stage_im_out(1409),
            product_re_out=>mul_re_out(1409),
            product_im_out=>mul_im_out(1409)
        );

    UMUL_1410 : complex_multiplier
    generic map(
            re_multiplicator=>15790, --- 0.963745117188 + j-0.266662597656
            im_multiplicator=>-4369
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1410),
            data_im_in=>first_stage_im_out(1410),
            product_re_out=>mul_re_out(1410),
            product_im_out=>mul_im_out(1410)
        );

    UMUL_1411 : complex_multiplier
    generic map(
            re_multiplicator=>15058, --- 0.919067382812 + j-0.393981933594
            im_multiplicator=>-6455
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1411),
            data_im_in=>first_stage_im_out(1411),
            product_re_out=>mul_re_out(1411),
            product_im_out=>mul_im_out(1411)
        );

    UMUL_1412 : complex_multiplier
    generic map(
            re_multiplicator=>14053, --- 0.857727050781 + j-0.514099121094
            im_multiplicator=>-8423
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1412),
            data_im_in=>first_stage_im_out(1412),
            product_re_out=>mul_re_out(1412),
            product_im_out=>mul_im_out(1412)
        );

    UMUL_1413 : complex_multiplier
    generic map(
            re_multiplicator=>12791, --- 0.780700683594 + j-0.624816894531
            im_multiplicator=>-10237
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1413),
            data_im_in=>first_stage_im_out(1413),
            product_re_out=>mul_re_out(1413),
            product_im_out=>mul_im_out(1413)
        );

    UMUL_1414 : complex_multiplier
    generic map(
            re_multiplicator=>11297, --- 0.689514160156 + j-0.724243164062
            im_multiplicator=>-11866
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1414),
            data_im_in=>first_stage_im_out(1414),
            product_re_out=>mul_re_out(1414),
            product_im_out=>mul_im_out(1414)
        );

    UMUL_1415 : complex_multiplier
    generic map(
            re_multiplicator=>9597, --- 0.585754394531 + j-0.810424804688
            im_multiplicator=>-13278
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1415),
            data_im_in=>first_stage_im_out(1415),
            product_re_out=>mul_re_out(1415),
            product_im_out=>mul_im_out(1415)
        );

    UMUL_1416 : complex_multiplier
    generic map(
            re_multiplicator=>7723, --- 0.471374511719 + j-0.881896972656
            im_multiplicator=>-14449
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1416),
            data_im_in=>first_stage_im_out(1416),
            product_re_out=>mul_re_out(1416),
            product_im_out=>mul_im_out(1416)
        );

    UMUL_1417 : complex_multiplier
    generic map(
            re_multiplicator=>5708, --- 0.348388671875 + j-0.937316894531
            im_multiplicator=>-15357
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1417),
            data_im_in=>first_stage_im_out(1417),
            product_re_out=>mul_re_out(1417),
            product_im_out=>mul_im_out(1417)
        );

    UMUL_1418 : complex_multiplier
    generic map(
            re_multiplicator=>3589, --- 0.219055175781 + j-0.975646972656
            im_multiplicator=>-15985
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1418),
            data_im_in=>first_stage_im_out(1418),
            product_re_out=>mul_re_out(1418),
            product_im_out=>mul_im_out(1418)
        );

    UMUL_1419 : complex_multiplier
    generic map(
            re_multiplicator=>1405, --- 0.0857543945312 + j-0.996276855469
            im_multiplicator=>-16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1419),
            data_im_in=>first_stage_im_out(1419),
            product_re_out=>mul_re_out(1419),
            product_im_out=>mul_im_out(1419)
        );

    UMUL_1420 : complex_multiplier
    generic map(
            re_multiplicator=>-803, --- -0.0490112304688 + j-0.998779296875
            im_multiplicator=>-16364
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1420),
            data_im_in=>first_stage_im_out(1420),
            product_re_out=>mul_re_out(1420),
            product_im_out=>mul_im_out(1420)
        );

    UMUL_1421 : complex_multiplier
    generic map(
            re_multiplicator=>-2998, --- -0.182983398438 + j-0.983093261719
            im_multiplicator=>-16107
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1421),
            data_im_in=>first_stage_im_out(1421),
            product_re_out=>mul_re_out(1421),
            product_im_out=>mul_im_out(1421)
        );

    UMUL_1422 : complex_multiplier
    generic map(
            re_multiplicator=>-5139, --- -0.313659667969 + j-0.949523925781
            im_multiplicator=>-15557
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1422),
            data_im_in=>first_stage_im_out(1422),
            product_re_out=>mul_re_out(1422),
            product_im_out=>mul_im_out(1422)
        );

    UMUL_1423 : complex_multiplier
    generic map(
            re_multiplicator=>-7186, --- -0.438598632812 + j-0.898620605469
            im_multiplicator=>-14723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1423),
            data_im_in=>first_stage_im_out(1423),
            product_re_out=>mul_re_out(1423),
            product_im_out=>mul_im_out(1423)
        );

    UMUL_1424 : complex_multiplier
    generic map(
            re_multiplicator=>-9102, --- -0.555541992188 + j-0.831420898438
            im_multiplicator=>-13622
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1424),
            data_im_in=>first_stage_im_out(1424),
            product_re_out=>mul_re_out(1424),
            product_im_out=>mul_im_out(1424)
        );

    UMUL_1425 : complex_multiplier
    generic map(
            re_multiplicator=>-10853, --- -0.662414550781 + j-0.749084472656
            im_multiplicator=>-12273
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1425),
            data_im_in=>first_stage_im_out(1425),
            product_re_out=>mul_re_out(1425),
            product_im_out=>mul_im_out(1425)
        );

    UMUL_1426 : complex_multiplier
    generic map(
            re_multiplicator=>-12406, --- -0.757202148438 + j-0.653137207031
            im_multiplicator=>-10701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1426),
            data_im_in=>first_stage_im_out(1426),
            product_re_out=>mul_re_out(1426),
            product_im_out=>mul_im_out(1426)
        );

    UMUL_1427 : complex_multiplier
    generic map(
            re_multiplicator=>-13733, --- -0.838195800781 + j-0.545288085938
            im_multiplicator=>-8934
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1427),
            data_im_in=>first_stage_im_out(1427),
            product_re_out=>mul_re_out(1427),
            product_im_out=>mul_im_out(1427)
        );

    UMUL_1428 : complex_multiplier
    generic map(
            re_multiplicator=>-14810, --- -0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1428),
            data_im_in=>first_stage_im_out(1428),
            product_re_out=>mul_re_out(1428),
            product_im_out=>mul_im_out(1428)
        );

    UMUL_1429 : complex_multiplier
    generic map(
            re_multiplicator=>-15618, --- -0.953247070312 + j-0.302001953125
            im_multiplicator=>-4948
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1429),
            data_im_in=>first_stage_im_out(1429),
            product_re_out=>mul_re_out(1429),
            product_im_out=>mul_im_out(1429)
        );

    UMUL_1430 : complex_multiplier
    generic map(
            re_multiplicator=>-16142, --- -0.985229492188 + j-0.170959472656
            im_multiplicator=>-2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1430),
            data_im_in=>first_stage_im_out(1430),
            product_re_out=>mul_re_out(1430),
            product_im_out=>mul_im_out(1430)
        );

    UMUL_1431 : complex_multiplier
    generic map(
            re_multiplicator=>-16372, --- -0.999267578125 + j-0.0368041992188
            im_multiplicator=>-603
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1431),
            data_im_in=>first_stage_im_out(1431),
            product_re_out=>mul_re_out(1431),
            product_im_out=>mul_im_out(1431)
        );

    UMUL_1432 : complex_multiplier
    generic map(
            re_multiplicator=>-16305, --- -0.995178222656 + j0.0979614257812
            im_multiplicator=>1605
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1432),
            data_im_in=>first_stage_im_out(1432),
            product_re_out=>mul_re_out(1432),
            product_im_out=>mul_im_out(1432)
        );

    UMUL_1433 : complex_multiplier
    generic map(
            re_multiplicator=>-15940, --- -0.972900390625 + j0.231018066406
            im_multiplicator=>3785
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1433),
            data_im_in=>first_stage_im_out(1433),
            product_re_out=>mul_re_out(1433),
            product_im_out=>mul_im_out(1433)
        );

    UMUL_1434 : complex_multiplier
    generic map(
            re_multiplicator=>-15286, --- -0.932983398438 + j0.35986328125
            im_multiplicator=>5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1434),
            data_im_in=>first_stage_im_out(1434),
            product_re_out=>mul_re_out(1434),
            product_im_out=>mul_im_out(1434)
        );

    UMUL_1435 : complex_multiplier
    generic map(
            re_multiplicator=>-14353, --- -0.876037597656 + j0.482177734375
            im_multiplicator=>7900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1435),
            data_im_in=>first_stage_im_out(1435),
            product_re_out=>mul_re_out(1435),
            product_im_out=>mul_im_out(1435)
        );

    UMUL_1436 : complex_multiplier
    generic map(
            re_multiplicator=>-13159, --- -0.803161621094 + j0.595642089844
            im_multiplicator=>9759
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1436),
            data_im_in=>first_stage_im_out(1436),
            product_re_out=>mul_re_out(1436),
            product_im_out=>mul_im_out(1436)
        );

    UMUL_1437 : complex_multiplier
    generic map(
            re_multiplicator=>-11726, --- -0.715698242188 + j0.698364257812
            im_multiplicator=>11442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1437),
            data_im_in=>first_stage_im_out(1437),
            product_re_out=>mul_re_out(1437),
            product_im_out=>mul_im_out(1437)
        );

    UMUL_1438 : complex_multiplier
    generic map(
            re_multiplicator=>-10079, --- -0.615173339844 + j0.788330078125
            im_multiplicator=>12916
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1438),
            data_im_in=>first_stage_im_out(1438),
            product_re_out=>mul_re_out(1438),
            product_im_out=>mul_im_out(1438)
        );

    UMUL_1439 : complex_multiplier
    generic map(
            re_multiplicator=>-8249, --- -0.503479003906 + j0.863952636719
            im_multiplicator=>14155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1439),
            data_im_in=>first_stage_im_out(1439),
            product_re_out=>mul_re_out(1439),
            product_im_out=>mul_im_out(1439)
        );

    UDELAY_1440_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1440),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1440)
        );
    UDELAY_1440_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1440),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1440)
        );
    USHIFTER_1440_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1440),
            data_out=>mul_re_out(1440)
        );
    USHIFTER_1440_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1440),
            data_out=>mul_im_out(1440)
        );

    UMUL_1441 : complex_multiplier
    generic map(
            re_multiplicator=>16228, --- 0.990478515625 + j-0.137573242188
            im_multiplicator=>-2254
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1441),
            data_im_in=>first_stage_im_out(1441),
            product_re_out=>mul_re_out(1441),
            product_im_out=>mul_im_out(1441)
        );

    UMUL_1442 : complex_multiplier
    generic map(
            re_multiplicator=>15763, --- 0.962097167969 + j-0.272583007812
            im_multiplicator=>-4466
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1442),
            data_im_in=>first_stage_im_out(1442),
            product_re_out=>mul_re_out(1442),
            product_im_out=>mul_im_out(1442)
        );

    UMUL_1443 : complex_multiplier
    generic map(
            re_multiplicator=>14998, --- 0.915405273438 + j-0.402404785156
            im_multiplicator=>-6593
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1443),
            data_im_in=>first_stage_im_out(1443),
            product_re_out=>mul_re_out(1443),
            product_im_out=>mul_im_out(1443)
        );

    UMUL_1444 : complex_multiplier
    generic map(
            re_multiplicator=>13948, --- 0.851318359375 + j-0.524536132812
            im_multiplicator=>-8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1444),
            data_im_in=>first_stage_im_out(1444),
            product_re_out=>mul_re_out(1444),
            product_im_out=>mul_im_out(1444)
        );

    UMUL_1445 : complex_multiplier
    generic map(
            re_multiplicator=>12633, --- 0.771057128906 + j-0.63671875
            im_multiplicator=>-10432
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1445),
            data_im_in=>first_stage_im_out(1445),
            product_re_out=>mul_re_out(1445),
            product_im_out=>mul_im_out(1445)
        );

    UMUL_1446 : complex_multiplier
    generic map(
            re_multiplicator=>11077, --- 0.676086425781 + j-0.73681640625
            im_multiplicator=>-12072
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1446),
            data_im_in=>first_stage_im_out(1446),
            product_re_out=>mul_re_out(1446),
            product_im_out=>mul_im_out(1446)
        );

    UMUL_1447 : complex_multiplier
    generic map(
            re_multiplicator=>9310, --- 0.568237304688 + j-0.822814941406
            im_multiplicator=>-13481
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1447),
            data_im_in=>first_stage_im_out(1447),
            product_re_out=>mul_re_out(1447),
            product_im_out=>mul_im_out(1447)
        );

    UMUL_1448 : complex_multiplier
    generic map(
            re_multiplicator=>7366, --- 0.449584960938 + j-0.893188476562
            im_multiplicator=>-14634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1448),
            data_im_in=>first_stage_im_out(1448),
            product_re_out=>mul_re_out(1448),
            product_im_out=>mul_im_out(1448)
        );

    UMUL_1449 : complex_multiplier
    generic map(
            re_multiplicator=>5282, --- 0.322387695312 + j-0.946594238281
            im_multiplicator=>-15509
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1449),
            data_im_in=>first_stage_im_out(1449),
            product_re_out=>mul_re_out(1449),
            product_im_out=>mul_im_out(1449)
        );

    UMUL_1450 : complex_multiplier
    generic map(
            re_multiplicator=>3097, --- 0.189025878906 + j-0.98193359375
            im_multiplicator=>-16088
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1450),
            data_im_in=>first_stage_im_out(1450),
            product_re_out=>mul_re_out(1450),
            product_im_out=>mul_im_out(1450)
        );

    UMUL_1451 : complex_multiplier
    generic map(
            re_multiplicator=>854, --- 0.0521240234375 + j-0.998596191406
            im_multiplicator=>-16361
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1451),
            data_im_in=>first_stage_im_out(1451),
            product_re_out=>mul_re_out(1451),
            product_im_out=>mul_im_out(1451)
        );

    UMUL_1452 : complex_multiplier
    generic map(
            re_multiplicator=>-1405, --- -0.0857543945312 + j-0.996276855469
            im_multiplicator=>-16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1452),
            data_im_in=>first_stage_im_out(1452),
            product_re_out=>mul_re_out(1452),
            product_im_out=>mul_im_out(1452)
        );

    UMUL_1453 : complex_multiplier
    generic map(
            re_multiplicator=>-3638, --- -0.222045898438 + j-0.974975585938
            im_multiplicator=>-15974
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1453),
            data_im_in=>first_stage_im_out(1453),
            product_re_out=>mul_re_out(1453),
            product_im_out=>mul_im_out(1453)
        );

    UMUL_1454 : complex_multiplier
    generic map(
            re_multiplicator=>-5802, --- -0.354125976562 + j-0.935180664062
            im_multiplicator=>-15322
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1454),
            data_im_in=>first_stage_im_out(1454),
            product_re_out=>mul_re_out(1454),
            product_im_out=>mul_im_out(1454)
        );

    UMUL_1455 : complex_multiplier
    generic map(
            re_multiplicator=>-7856, --- -0.4794921875 + j-0.877502441406
            im_multiplicator=>-14377
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1455),
            data_im_in=>first_stage_im_out(1455),
            product_re_out=>mul_re_out(1455),
            product_im_out=>mul_im_out(1455)
        );

    UMUL_1456 : complex_multiplier
    generic map(
            re_multiplicator=>-9759, --- -0.595642089844 + j-0.803161621094
            im_multiplicator=>-13159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1456),
            data_im_in=>first_stage_im_out(1456),
            product_re_out=>mul_re_out(1456),
            product_im_out=>mul_im_out(1456)
        );

    UMUL_1457 : complex_multiplier
    generic map(
            re_multiplicator=>-11478, --- -0.700561523438 + j-0.713562011719
            im_multiplicator=>-11691
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1457),
            data_im_in=>first_stage_im_out(1457),
            product_re_out=>mul_re_out(1457),
            product_im_out=>mul_im_out(1457)
        );

    UMUL_1458 : complex_multiplier
    generic map(
            re_multiplicator=>-12977, --- -0.792053222656 + j-0.6103515625
            im_multiplicator=>-10000
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1458),
            data_im_in=>first_stage_im_out(1458),
            product_re_out=>mul_re_out(1458),
            product_im_out=>mul_im_out(1458)
        );

    UMUL_1459 : complex_multiplier
    generic map(
            re_multiplicator=>-14230, --- -0.868530273438 + j-0.495544433594
            im_multiplicator=>-8119
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1459),
            data_im_in=>first_stage_im_out(1459),
            product_re_out=>mul_re_out(1459),
            product_im_out=>mul_im_out(1459)
        );

    UMUL_1460 : complex_multiplier
    generic map(
            re_multiplicator=>-15212, --- -0.928466796875 + j-0.371276855469
            im_multiplicator=>-6083
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1460),
            data_im_in=>first_stage_im_out(1460),
            product_re_out=>mul_re_out(1460),
            product_im_out=>mul_im_out(1460)
        );

    UMUL_1461 : complex_multiplier
    generic map(
            re_multiplicator=>-15905, --- -0.970764160156 + j-0.239990234375
            im_multiplicator=>-3932
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1461),
            data_im_in=>first_stage_im_out(1461),
            product_re_out=>mul_re_out(1461),
            product_im_out=>mul_im_out(1461)
        );

    UMUL_1462 : complex_multiplier
    generic map(
            re_multiplicator=>-16294, --- -0.994506835938 + j-0.104064941406
            im_multiplicator=>-1705
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1462),
            data_im_in=>first_stage_im_out(1462),
            product_re_out=>mul_re_out(1462),
            product_im_out=>mul_im_out(1462)
        );

    UMUL_1463 : complex_multiplier
    generic map(
            re_multiplicator=>-16374, --- -0.999389648438 + j0.03369140625
            im_multiplicator=>552
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1463),
            data_im_in=>first_stage_im_out(1463),
            product_re_out=>mul_re_out(1463),
            product_im_out=>mul_im_out(1463)
        );

    UMUL_1464 : complex_multiplier
    generic map(
            re_multiplicator=>-16142, --- -0.985229492188 + j0.170959472656
            im_multiplicator=>2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1464),
            data_im_in=>first_stage_im_out(1464),
            product_re_out=>mul_re_out(1464),
            product_im_out=>mul_im_out(1464)
        );

    UMUL_1465 : complex_multiplier
    generic map(
            re_multiplicator=>-15603, --- -0.952331542969 + j0.304870605469
            im_multiplicator=>4995
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1465),
            data_im_in=>first_stage_im_out(1465),
            product_re_out=>mul_re_out(1465),
            product_im_out=>mul_im_out(1465)
        );

    UMUL_1466 : complex_multiplier
    generic map(
            re_multiplicator=>-14767, --- -0.901306152344 + j0.433044433594
            im_multiplicator=>7095
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1466),
            data_im_in=>first_stage_im_out(1466),
            product_re_out=>mul_re_out(1466),
            product_im_out=>mul_im_out(1466)
        );

    UMUL_1467 : complex_multiplier
    generic map(
            re_multiplicator=>-13650, --- -0.833129882812 + j0.552978515625
            im_multiplicator=>9060
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1467),
            data_im_in=>first_stage_im_out(1467),
            product_re_out=>mul_re_out(1467),
            product_im_out=>mul_im_out(1467)
        );

    UMUL_1468 : complex_multiplier
    generic map(
            re_multiplicator=>-12273, --- -0.749084472656 + j0.662414550781
            im_multiplicator=>10853
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1468),
            data_im_in=>first_stage_im_out(1468),
            product_re_out=>mul_re_out(1468),
            product_im_out=>mul_im_out(1468)
        );

    UMUL_1469 : complex_multiplier
    generic map(
            re_multiplicator=>-10663, --- -0.650817871094 + j0.759155273438
            im_multiplicator=>12438
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1469),
            data_im_in=>first_stage_im_out(1469),
            product_re_out=>mul_re_out(1469),
            product_im_out=>mul_im_out(1469)
        );

    UMUL_1470 : complex_multiplier
    generic map(
            re_multiplicator=>-8850, --- -0.540161132812 + j0.841552734375
            im_multiplicator=>13788
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1470),
            data_im_in=>first_stage_im_out(1470),
            product_re_out=>mul_re_out(1470),
            product_im_out=>mul_im_out(1470)
        );

    UMUL_1471 : complex_multiplier
    generic map(
            re_multiplicator=>-6868, --- -0.419189453125 + j0.907836914062
            im_multiplicator=>14874
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1471),
            data_im_in=>first_stage_im_out(1471),
            product_re_out=>mul_re_out(1471),
            product_im_out=>mul_im_out(1471)
        );

    UDELAY_1472_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1472),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1472)
        );
    UDELAY_1472_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1472),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1472)
        );
    USHIFTER_1472_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1472),
            data_out=>mul_re_out(1472)
        );
    USHIFTER_1472_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1472),
            data_out=>mul_im_out(1472)
        );

    UMUL_1473 : complex_multiplier
    generic map(
            re_multiplicator=>16221, --- 0.990051269531 + j-0.140625
            im_multiplicator=>-2304
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1473),
            data_im_in=>first_stage_im_out(1473),
            product_re_out=>mul_re_out(1473),
            product_im_out=>mul_im_out(1473)
        );

    UMUL_1474 : complex_multiplier
    generic map(
            re_multiplicator=>15735, --- 0.960388183594 + j-0.278503417969
            im_multiplicator=>-4563
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1474),
            data_im_in=>first_stage_im_out(1474),
            product_re_out=>mul_re_out(1474),
            product_im_out=>mul_im_out(1474)
        );

    UMUL_1475 : complex_multiplier
    generic map(
            re_multiplicator=>14937, --- 0.911682128906 + j-0.410827636719
            im_multiplicator=>-6731
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1475),
            data_im_in=>first_stage_im_out(1475),
            product_re_out=>mul_re_out(1475),
            product_im_out=>mul_im_out(1475)
        );

    UMUL_1476 : complex_multiplier
    generic map(
            re_multiplicator=>13842, --- 0.844848632812 + j-0.534973144531
            im_multiplicator=>-8765
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1476),
            data_im_in=>first_stage_im_out(1476),
            product_re_out=>mul_re_out(1476),
            product_im_out=>mul_im_out(1476)
        );

    UMUL_1477 : complex_multiplier
    generic map(
            re_multiplicator=>12471, --- 0.761169433594 + j-0.648498535156
            im_multiplicator=>-10625
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1477),
            data_im_in=>first_stage_im_out(1477),
            product_re_out=>mul_re_out(1477),
            product_im_out=>mul_im_out(1477)
        );

    UMUL_1478 : complex_multiplier
    generic map(
            re_multiplicator=>10853, --- 0.662414550781 + j-0.749084472656
            im_multiplicator=>-12273
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1478),
            data_im_in=>first_stage_im_out(1478),
            product_re_out=>mul_re_out(1478),
            product_im_out=>mul_im_out(1478)
        );

    UMUL_1479 : complex_multiplier
    generic map(
            re_multiplicator=>9018, --- 0.550415039062 + j-0.834838867188
            im_multiplicator=>-13678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1479),
            data_im_in=>first_stage_im_out(1479),
            product_re_out=>mul_re_out(1479),
            product_im_out=>mul_im_out(1479)
        );

    UMUL_1480 : complex_multiplier
    generic map(
            re_multiplicator=>7005, --- 0.427551269531 + j-0.903930664062
            im_multiplicator=>-14810
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1480),
            data_im_in=>first_stage_im_out(1480),
            product_re_out=>mul_re_out(1480),
            product_im_out=>mul_im_out(1480)
        );

    UMUL_1481 : complex_multiplier
    generic map(
            re_multiplicator=>4852, --- 0.296142578125 + j-0.955139160156
            im_multiplicator=>-15649
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1481),
            data_im_in=>first_stage_im_out(1481),
            product_re_out=>mul_re_out(1481),
            product_im_out=>mul_im_out(1481)
        );

    UMUL_1482 : complex_multiplier
    generic map(
            re_multiplicator=>2602, --- 0.158813476562 + j-0.987243652344
            im_multiplicator=>-16175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1482),
            data_im_in=>first_stage_im_out(1482),
            product_re_out=>mul_re_out(1482),
            product_im_out=>mul_im_out(1482)
        );

    UMUL_1483 : complex_multiplier
    generic map(
            re_multiplicator=>301, --- 0.0183715820312 + j-0.999816894531
            im_multiplicator=>-16381
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1483),
            data_im_in=>first_stage_im_out(1483),
            product_re_out=>mul_re_out(1483),
            product_im_out=>mul_im_out(1483)
        );

    UMUL_1484 : complex_multiplier
    generic map(
            re_multiplicator=>-2005, --- -0.122375488281 + j-0.992431640625
            im_multiplicator=>-16260
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1484),
            data_im_in=>first_stage_im_out(1484),
            product_re_out=>mul_re_out(1484),
            product_im_out=>mul_im_out(1484)
        );

    UMUL_1485 : complex_multiplier
    generic map(
            re_multiplicator=>-4272, --- -0.2607421875 + j-0.965393066406
            im_multiplicator=>-15817
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1485),
            data_im_in=>first_stage_im_out(1485),
            product_re_out=>mul_re_out(1485),
            product_im_out=>mul_im_out(1485)
        );

    UMUL_1486 : complex_multiplier
    generic map(
            re_multiplicator=>-6455, --- -0.393981933594 + j-0.919067382812
            im_multiplicator=>-15058
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1486),
            data_im_in=>first_stage_im_out(1486),
            product_re_out=>mul_re_out(1486),
            product_im_out=>mul_im_out(1486)
        );

    UMUL_1487 : complex_multiplier
    generic map(
            re_multiplicator=>-8509, --- -0.519348144531 + j-0.854553222656
            im_multiplicator=>-14001
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1487),
            data_im_in=>first_stage_im_out(1487),
            product_re_out=>mul_re_out(1487),
            product_im_out=>mul_im_out(1487)
        );

    UMUL_1488 : complex_multiplier
    generic map(
            re_multiplicator=>-10393, --- -0.634338378906 + j-0.773010253906
            im_multiplicator=>-12665
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1488),
            data_im_in=>first_stage_im_out(1488),
            product_re_out=>mul_re_out(1488),
            product_im_out=>mul_im_out(1488)
        );

    UMUL_1489 : complex_multiplier
    generic map(
            re_multiplicator=>-12072, --- -0.73681640625 + j-0.676086425781
            im_multiplicator=>-11077
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1489),
            data_im_in=>first_stage_im_out(1489),
            product_re_out=>mul_re_out(1489),
            product_im_out=>mul_im_out(1489)
        );

    UMUL_1490 : complex_multiplier
    generic map(
            re_multiplicator=>-13510, --- -0.824584960938 + j-0.565673828125
            im_multiplicator=>-9268
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1490),
            data_im_in=>first_stage_im_out(1490),
            product_re_out=>mul_re_out(1490),
            product_im_out=>mul_im_out(1490)
        );

    UMUL_1491 : complex_multiplier
    generic map(
            re_multiplicator=>-14679, --- -0.895935058594 + j-0.444091796875
            im_multiplicator=>-7276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1491),
            data_im_in=>first_stage_im_out(1491),
            product_re_out=>mul_re_out(1491),
            product_im_out=>mul_im_out(1491)
        );

    UMUL_1492 : complex_multiplier
    generic map(
            re_multiplicator=>-15557, --- -0.949523925781 + j-0.313659667969
            im_multiplicator=>-5139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1492),
            data_im_in=>first_stage_im_out(1492),
            product_re_out=>mul_re_out(1492),
            product_im_out=>mul_im_out(1492)
        );

    UMUL_1493 : complex_multiplier
    generic map(
            re_multiplicator=>-16125, --- -0.984191894531 + j-0.177001953125
            im_multiplicator=>-2900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1493),
            data_im_in=>first_stage_im_out(1493),
            product_re_out=>mul_re_out(1493),
            product_im_out=>mul_im_out(1493)
        );

    UMUL_1494 : complex_multiplier
    generic map(
            re_multiplicator=>-16372, --- -0.999267578125 + j-0.0368041992188
            im_multiplicator=>-603
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1494),
            data_im_in=>first_stage_im_out(1494),
            product_re_out=>mul_re_out(1494),
            product_im_out=>mul_im_out(1494)
        );

    UMUL_1495 : complex_multiplier
    generic map(
            re_multiplicator=>-16294, --- -0.994506835938 + j0.104064941406
            im_multiplicator=>1705
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1495),
            data_im_in=>first_stage_im_out(1495),
            product_re_out=>mul_re_out(1495),
            product_im_out=>mul_im_out(1495)
        );

    UMUL_1496 : complex_multiplier
    generic map(
            re_multiplicator=>-15892, --- -0.969970703125 + j0.242919921875
            im_multiplicator=>3980
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1496),
            data_im_in=>first_stage_im_out(1496),
            product_re_out=>mul_re_out(1496),
            product_im_out=>mul_im_out(1496)
        );

    UMUL_1497 : complex_multiplier
    generic map(
            re_multiplicator=>-15175, --- -0.926208496094 + j0.376953125
            im_multiplicator=>6176
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1497),
            data_im_in=>first_stage_im_out(1497),
            product_re_out=>mul_re_out(1497),
            product_im_out=>mul_im_out(1497)
        );

    UMUL_1498 : complex_multiplier
    generic map(
            re_multiplicator=>-14155, --- -0.863952636719 + j0.503479003906
            im_multiplicator=>8249
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1498),
            data_im_in=>first_stage_im_out(1498),
            product_re_out=>mul_re_out(1498),
            product_im_out=>mul_im_out(1498)
        );

    UMUL_1499 : complex_multiplier
    generic map(
            re_multiplicator=>-12854, --- -0.784545898438 + j0.620056152344
            im_multiplicator=>10159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1499),
            data_im_in=>first_stage_im_out(1499),
            product_re_out=>mul_re_out(1499),
            product_im_out=>mul_im_out(1499)
        );

    UMUL_1500 : complex_multiplier
    generic map(
            re_multiplicator=>-11297, --- -0.689514160156 + j0.724243164062
            im_multiplicator=>11866
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1500),
            data_im_in=>first_stage_im_out(1500),
            product_re_out=>mul_re_out(1500),
            product_im_out=>mul_im_out(1500)
        );

    UMUL_1501 : complex_multiplier
    generic map(
            re_multiplicator=>-9516, --- -0.580810546875 + j0.814025878906
            im_multiplicator=>13337
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1501),
            data_im_in=>first_stage_im_out(1501),
            product_re_out=>mul_re_out(1501),
            product_im_out=>mul_im_out(1501)
        );

    UMUL_1502 : complex_multiplier
    generic map(
            re_multiplicator=>-7545, --- -0.460510253906 + j0.887634277344
            im_multiplicator=>14543
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1502),
            data_im_in=>first_stage_im_out(1502),
            product_re_out=>mul_re_out(1502),
            product_im_out=>mul_im_out(1502)
        );

    UMUL_1503 : complex_multiplier
    generic map(
            re_multiplicator=>-5424, --- -0.3310546875 + j0.943542480469
            im_multiplicator=>15459
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1503),
            data_im_in=>first_stage_im_out(1503),
            product_re_out=>mul_re_out(1503),
            product_im_out=>mul_im_out(1503)
        );

    UDELAY_1504_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1504),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1504)
        );
    UDELAY_1504_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1504),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1504)
        );
    USHIFTER_1504_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1504),
            data_out=>mul_re_out(1504)
        );
    USHIFTER_1504_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1504),
            data_out=>mul_im_out(1504)
        );

    UMUL_1505 : complex_multiplier
    generic map(
            re_multiplicator=>16213, --- 0.989562988281 + j-0.143676757812
            im_multiplicator=>-2354
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1505),
            data_im_in=>first_stage_im_out(1505),
            product_re_out=>mul_re_out(1505),
            product_im_out=>mul_im_out(1505)
        );

    UMUL_1506 : complex_multiplier
    generic map(
            re_multiplicator=>15707, --- 0.958679199219 + j-0.284362792969
            im_multiplicator=>-4659
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1506),
            data_im_in=>first_stage_im_out(1506),
            product_re_out=>mul_re_out(1506),
            product_im_out=>mul_im_out(1506)
        );

    UMUL_1507 : complex_multiplier
    generic map(
            re_multiplicator=>14874, --- 0.907836914062 + j-0.419189453125
            im_multiplicator=>-6868
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1507),
            data_im_in=>first_stage_im_out(1507),
            product_re_out=>mul_re_out(1507),
            product_im_out=>mul_im_out(1507)
        );

    UMUL_1508 : complex_multiplier
    generic map(
            re_multiplicator=>13733, --- 0.838195800781 + j-0.545288085938
            im_multiplicator=>-8934
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1508),
            data_im_in=>first_stage_im_out(1508),
            product_re_out=>mul_re_out(1508),
            product_im_out=>mul_im_out(1508)
        );

    UMUL_1509 : complex_multiplier
    generic map(
            re_multiplicator=>12307, --- 0.751159667969 + j-0.660095214844
            im_multiplicator=>-10815
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1509),
            data_im_in=>first_stage_im_out(1509),
            product_re_out=>mul_re_out(1509),
            product_im_out=>mul_im_out(1509)
        );

    UMUL_1510 : complex_multiplier
    generic map(
            re_multiplicator=>10625, --- 0.648498535156 + j-0.761169433594
            im_multiplicator=>-12471
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1510),
            data_im_in=>first_stage_im_out(1510),
            product_re_out=>mul_re_out(1510),
            product_im_out=>mul_im_out(1510)
        );

    UMUL_1511 : complex_multiplier
    generic map(
            re_multiplicator=>8722, --- 0.532348632812 + j-0.846435546875
            im_multiplicator=>-13868
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1511),
            data_im_in=>first_stage_im_out(1511),
            product_re_out=>mul_re_out(1511),
            product_im_out=>mul_im_out(1511)
        );

    UMUL_1512 : complex_multiplier
    generic map(
            re_multiplicator=>6639, --- 0.405212402344 + j-0.914184570312
            im_multiplicator=>-14978
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1512),
            data_im_in=>first_stage_im_out(1512),
            product_re_out=>mul_re_out(1512),
            product_im_out=>mul_im_out(1512)
        );

    UMUL_1513 : complex_multiplier
    generic map(
            re_multiplicator=>4418, --- 0.269653320312 + j-0.962951660156
            im_multiplicator=>-15777
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1513),
            data_im_in=>first_stage_im_out(1513),
            product_re_out=>mul_re_out(1513),
            product_im_out=>mul_im_out(1513)
        );

    UMUL_1514 : complex_multiplier
    generic map(
            re_multiplicator=>2105, --- 0.128479003906 + j-0.99169921875
            im_multiplicator=>-16248
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1514),
            data_im_in=>first_stage_im_out(1514),
            product_re_out=>mul_re_out(1514),
            product_im_out=>mul_im_out(1514)
        );

    UMUL_1515 : complex_multiplier
    generic map(
            re_multiplicator=>-251, --- -0.0153198242188 + j-0.999877929688
            im_multiplicator=>-16382
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1515),
            data_im_in=>first_stage_im_out(1515),
            product_re_out=>mul_re_out(1515),
            product_im_out=>mul_im_out(1515)
        );

    UMUL_1516 : complex_multiplier
    generic map(
            re_multiplicator=>-2602, --- -0.158813476562 + j-0.987243652344
            im_multiplicator=>-16175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1516),
            data_im_in=>first_stage_im_out(1516),
            product_re_out=>mul_re_out(1516),
            product_im_out=>mul_im_out(1516)
        );

    UMUL_1517 : complex_multiplier
    generic map(
            re_multiplicator=>-4900, --- -0.299072265625 + j-0.954223632812
            im_multiplicator=>-15634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1517),
            data_im_in=>first_stage_im_out(1517),
            product_re_out=>mul_re_out(1517),
            product_im_out=>mul_im_out(1517)
        );

    UMUL_1518 : complex_multiplier
    generic map(
            re_multiplicator=>-7095, --- -0.433044433594 + j-0.901306152344
            im_multiplicator=>-14767
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1518),
            data_im_in=>first_stage_im_out(1518),
            product_re_out=>mul_re_out(1518),
            product_im_out=>mul_im_out(1518)
        );

    UMUL_1519 : complex_multiplier
    generic map(
            re_multiplicator=>-9144, --- -0.55810546875 + j-0.829711914062
            im_multiplicator=>-13594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1519),
            data_im_in=>first_stage_im_out(1519),
            product_re_out=>mul_re_out(1519),
            product_im_out=>mul_im_out(1519)
        );

    UMUL_1520 : complex_multiplier
    generic map(
            re_multiplicator=>-11002, --- -0.671508789062 + j-0.740905761719
            im_multiplicator=>-12139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1520),
            data_im_in=>first_stage_im_out(1520),
            product_re_out=>mul_re_out(1520),
            product_im_out=>mul_im_out(1520)
        );

    UMUL_1521 : complex_multiplier
    generic map(
            re_multiplicator=>-12633, --- -0.771057128906 + j-0.63671875
            im_multiplicator=>-10432
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1521),
            data_im_in=>first_stage_im_out(1521),
            product_re_out=>mul_re_out(1521),
            product_im_out=>mul_im_out(1521)
        );

    UMUL_1522 : complex_multiplier
    generic map(
            re_multiplicator=>-14001, --- -0.854553222656 + j-0.519348144531
            im_multiplicator=>-8509
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1522),
            data_im_in=>first_stage_im_out(1522),
            product_re_out=>mul_re_out(1522),
            product_im_out=>mul_im_out(1522)
        );

    UMUL_1523 : complex_multiplier
    generic map(
            re_multiplicator=>-15078, --- -0.920288085938 + j-0.39111328125
            im_multiplicator=>-6408
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1523),
            data_im_in=>first_stage_im_out(1523),
            product_re_out=>mul_re_out(1523),
            product_im_out=>mul_im_out(1523)
        );

    UMUL_1524 : complex_multiplier
    generic map(
            re_multiplicator=>-15842, --- -0.966918945312 + j-0.254821777344
            im_multiplicator=>-4175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1524),
            data_im_in=>first_stage_im_out(1524),
            product_re_out=>mul_re_out(1524),
            product_im_out=>mul_im_out(1524)
        );

    UMUL_1525 : complex_multiplier
    generic map(
            re_multiplicator=>-16278, --- -0.993530273438 + j-0.113220214844
            im_multiplicator=>-1855
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1525),
            data_im_in=>first_stage_im_out(1525),
            product_re_out=>mul_re_out(1525),
            product_im_out=>mul_im_out(1525)
        );

    UMUL_1526 : complex_multiplier
    generic map(
            re_multiplicator=>-16376, --- -0.99951171875 + j0.0306396484375
            im_multiplicator=>502
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1526),
            data_im_in=>first_stage_im_out(1526),
            product_re_out=>mul_re_out(1526),
            product_im_out=>mul_im_out(1526)
        );

    UMUL_1527 : complex_multiplier
    generic map(
            re_multiplicator=>-16134, --- -0.984741210938 + j0.173950195312
            im_multiplicator=>2850
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1527),
            data_im_in=>first_stage_im_out(1527),
            product_re_out=>mul_re_out(1527),
            product_im_out=>mul_im_out(1527)
        );

    UMUL_1528 : complex_multiplier
    generic map(
            re_multiplicator=>-15557, --- -0.949523925781 + j0.313659667969
            im_multiplicator=>5139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1528),
            data_im_in=>first_stage_im_out(1528),
            product_re_out=>mul_re_out(1528),
            product_im_out=>mul_im_out(1528)
        );

    UMUL_1529 : complex_multiplier
    generic map(
            re_multiplicator=>-14657, --- -0.894592285156 + j0.446838378906
            im_multiplicator=>7321
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1529),
            data_im_in=>first_stage_im_out(1529),
            product_re_out=>mul_re_out(1529),
            product_im_out=>mul_im_out(1529)
        );

    UMUL_1530 : complex_multiplier
    generic map(
            re_multiplicator=>-13452, --- -0.821044921875 + j0.570739746094
            im_multiplicator=>9351
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1530),
            data_im_in=>first_stage_im_out(1530),
            product_re_out=>mul_re_out(1530),
            product_im_out=>mul_im_out(1530)
        );

    UMUL_1531 : complex_multiplier
    generic map(
            re_multiplicator=>-11969, --- -0.730529785156 + j0.682800292969
            im_multiplicator=>11187
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1531),
            data_im_in=>first_stage_im_out(1531),
            product_re_out=>mul_re_out(1531),
            product_im_out=>mul_im_out(1531)
        );

    UMUL_1532 : complex_multiplier
    generic map(
            re_multiplicator=>-10237, --- -0.624816894531 + j0.780700683594
            im_multiplicator=>12791
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1532),
            data_im_in=>first_stage_im_out(1532),
            product_re_out=>mul_re_out(1532),
            product_im_out=>mul_im_out(1532)
        );

    UMUL_1533 : complex_multiplier
    generic map(
            re_multiplicator=>-8293, --- -0.506164550781 + j0.862365722656
            im_multiplicator=>14129
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1533),
            data_im_in=>first_stage_im_out(1533),
            product_re_out=>mul_re_out(1533),
            product_im_out=>mul_im_out(1533)
        );

    UMUL_1534 : complex_multiplier
    generic map(
            re_multiplicator=>-6176, --- -0.376953125 + j0.926208496094
            im_multiplicator=>15175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1534),
            data_im_in=>first_stage_im_out(1534),
            product_re_out=>mul_re_out(1534),
            product_im_out=>mul_im_out(1534)
        );

    UMUL_1535 : complex_multiplier
    generic map(
            re_multiplicator=>-3932, --- -0.239990234375 + j0.970764160156
            im_multiplicator=>15905
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1535),
            data_im_in=>first_stage_im_out(1535),
            product_re_out=>mul_re_out(1535),
            product_im_out=>mul_im_out(1535)
        );

    UDELAY_1536_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1536),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1536)
        );
    UDELAY_1536_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1536),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1536)
        );
    USHIFTER_1536_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1536),
            data_out=>mul_re_out(1536)
        );
    USHIFTER_1536_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1536),
            data_out=>mul_im_out(1536)
        );

    UMUL_1537 : complex_multiplier
    generic map(
            re_multiplicator=>16206, --- 0.989135742188 + j-0.146728515625
            im_multiplicator=>-2404
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1537),
            data_im_in=>first_stage_im_out(1537),
            product_re_out=>mul_re_out(1537),
            product_im_out=>mul_im_out(1537)
        );

    UMUL_1538 : complex_multiplier
    generic map(
            re_multiplicator=>15678, --- 0.956909179688 + j-0.290283203125
            im_multiplicator=>-4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1538),
            data_im_in=>first_stage_im_out(1538),
            product_re_out=>mul_re_out(1538),
            product_im_out=>mul_im_out(1538)
        );

    UMUL_1539 : complex_multiplier
    generic map(
            re_multiplicator=>14810, --- 0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1539),
            data_im_in=>first_stage_im_out(1539),
            product_re_out=>mul_re_out(1539),
            product_im_out=>mul_im_out(1539)
        );

    UMUL_1540 : complex_multiplier
    generic map(
            re_multiplicator=>13622, --- 0.831420898438 + j-0.555541992188
            im_multiplicator=>-9102
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1540),
            data_im_in=>first_stage_im_out(1540),
            product_re_out=>mul_re_out(1540),
            product_im_out=>mul_im_out(1540)
        );

    UMUL_1541 : complex_multiplier
    generic map(
            re_multiplicator=>12139, --- 0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1541),
            data_im_in=>first_stage_im_out(1541),
            product_re_out=>mul_re_out(1541),
            product_im_out=>mul_im_out(1541)
        );

    UMUL_1542 : complex_multiplier
    generic map(
            re_multiplicator=>10393, --- 0.634338378906 + j-0.773010253906
            im_multiplicator=>-12665
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1542),
            data_im_in=>first_stage_im_out(1542),
            product_re_out=>mul_re_out(1542),
            product_im_out=>mul_im_out(1542)
        );

    UMUL_1543 : complex_multiplier
    generic map(
            re_multiplicator=>8423, --- 0.514099121094 + j-0.857727050781
            im_multiplicator=>-14053
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1543),
            data_im_in=>first_stage_im_out(1543),
            product_re_out=>mul_re_out(1543),
            product_im_out=>mul_im_out(1543)
        );

    UMUL_1544 : complex_multiplier
    generic map(
            re_multiplicator=>6269, --- 0.382629394531 + j-0.923828125
            im_multiplicator=>-15136
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1544),
            data_im_in=>first_stage_im_out(1544),
            product_re_out=>mul_re_out(1544),
            product_im_out=>mul_im_out(1544)
        );

    UMUL_1545 : complex_multiplier
    generic map(
            re_multiplicator=>3980, --- 0.242919921875 + j-0.969970703125
            im_multiplicator=>-15892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1545),
            data_im_in=>first_stage_im_out(1545),
            product_re_out=>mul_re_out(1545),
            product_im_out=>mul_im_out(1545)
        );

    UMUL_1546 : complex_multiplier
    generic map(
            re_multiplicator=>1605, --- 0.0979614257812 + j-0.995178222656
            im_multiplicator=>-16305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1546),
            data_im_in=>first_stage_im_out(1546),
            product_re_out=>mul_re_out(1546),
            product_im_out=>mul_im_out(1546)
        );

    UMUL_1547 : complex_multiplier
    generic map(
            re_multiplicator=>-803, --- -0.0490112304688 + j-0.998779296875
            im_multiplicator=>-16364
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1547),
            data_im_in=>first_stage_im_out(1547),
            product_re_out=>mul_re_out(1547),
            product_im_out=>mul_im_out(1547)
        );

    UMUL_1548 : complex_multiplier
    generic map(
            re_multiplicator=>-3196, --- -0.195068359375 + j-0.980773925781
            im_multiplicator=>-16069
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1548),
            data_im_in=>first_stage_im_out(1548),
            product_re_out=>mul_re_out(1548),
            product_im_out=>mul_im_out(1548)
        );

    UMUL_1549 : complex_multiplier
    generic map(
            re_multiplicator=>-5519, --- -0.336853027344 + j-0.941528320312
            im_multiplicator=>-15426
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1549),
            data_im_in=>first_stage_im_out(1549),
            product_re_out=>mul_re_out(1549),
            product_im_out=>mul_im_out(1549)
        );

    UMUL_1550 : complex_multiplier
    generic map(
            re_multiplicator=>-7723, --- -0.471374511719 + j-0.881896972656
            im_multiplicator=>-14449
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1550),
            data_im_in=>first_stage_im_out(1550),
            product_re_out=>mul_re_out(1550),
            product_im_out=>mul_im_out(1550)
        );

    UMUL_1551 : complex_multiplier
    generic map(
            re_multiplicator=>-9759, --- -0.595642089844 + j-0.803161621094
            im_multiplicator=>-13159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1551),
            data_im_in=>first_stage_im_out(1551),
            product_re_out=>mul_re_out(1551),
            product_im_out=>mul_im_out(1551)
        );

    UMUL_1552 : complex_multiplier
    generic map(
            re_multiplicator=>-11585, --- -0.707092285156 + j-0.707092285156
            im_multiplicator=>-11585
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1552),
            data_im_in=>first_stage_im_out(1552),
            product_re_out=>mul_re_out(1552),
            product_im_out=>mul_im_out(1552)
        );

    UMUL_1553 : complex_multiplier
    generic map(
            re_multiplicator=>-13159, --- -0.803161621094 + j-0.595642089844
            im_multiplicator=>-9759
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1553),
            data_im_in=>first_stage_im_out(1553),
            product_re_out=>mul_re_out(1553),
            product_im_out=>mul_im_out(1553)
        );

    UMUL_1554 : complex_multiplier
    generic map(
            re_multiplicator=>-14449, --- -0.881896972656 + j-0.471374511719
            im_multiplicator=>-7723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1554),
            data_im_in=>first_stage_im_out(1554),
            product_re_out=>mul_re_out(1554),
            product_im_out=>mul_im_out(1554)
        );

    UMUL_1555 : complex_multiplier
    generic map(
            re_multiplicator=>-15426, --- -0.941528320312 + j-0.336853027344
            im_multiplicator=>-5519
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1555),
            data_im_in=>first_stage_im_out(1555),
            product_re_out=>mul_re_out(1555),
            product_im_out=>mul_im_out(1555)
        );

    UMUL_1556 : complex_multiplier
    generic map(
            re_multiplicator=>-16069, --- -0.980773925781 + j-0.195068359375
            im_multiplicator=>-3196
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1556),
            data_im_in=>first_stage_im_out(1556),
            product_re_out=>mul_re_out(1556),
            product_im_out=>mul_im_out(1556)
        );

    UMUL_1557 : complex_multiplier
    generic map(
            re_multiplicator=>-16364, --- -0.998779296875 + j-0.0490112304688
            im_multiplicator=>-803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1557),
            data_im_in=>first_stage_im_out(1557),
            product_re_out=>mul_re_out(1557),
            product_im_out=>mul_im_out(1557)
        );

    UMUL_1558 : complex_multiplier
    generic map(
            re_multiplicator=>-16305, --- -0.995178222656 + j0.0979614257812
            im_multiplicator=>1605
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1558),
            data_im_in=>first_stage_im_out(1558),
            product_re_out=>mul_re_out(1558),
            product_im_out=>mul_im_out(1558)
        );

    UMUL_1559 : complex_multiplier
    generic map(
            re_multiplicator=>-15892, --- -0.969970703125 + j0.242919921875
            im_multiplicator=>3980
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1559),
            data_im_in=>first_stage_im_out(1559),
            product_re_out=>mul_re_out(1559),
            product_im_out=>mul_im_out(1559)
        );

    UMUL_1560 : complex_multiplier
    generic map(
            re_multiplicator=>-15136, --- -0.923828125 + j0.382629394531
            im_multiplicator=>6269
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1560),
            data_im_in=>first_stage_im_out(1560),
            product_re_out=>mul_re_out(1560),
            product_im_out=>mul_im_out(1560)
        );

    UMUL_1561 : complex_multiplier
    generic map(
            re_multiplicator=>-14053, --- -0.857727050781 + j0.514099121094
            im_multiplicator=>8423
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1561),
            data_im_in=>first_stage_im_out(1561),
            product_re_out=>mul_re_out(1561),
            product_im_out=>mul_im_out(1561)
        );

    UMUL_1562 : complex_multiplier
    generic map(
            re_multiplicator=>-12665, --- -0.773010253906 + j0.634338378906
            im_multiplicator=>10393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1562),
            data_im_in=>first_stage_im_out(1562),
            product_re_out=>mul_re_out(1562),
            product_im_out=>mul_im_out(1562)
        );

    UMUL_1563 : complex_multiplier
    generic map(
            re_multiplicator=>-11002, --- -0.671508789062 + j0.740905761719
            im_multiplicator=>12139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1563),
            data_im_in=>first_stage_im_out(1563),
            product_re_out=>mul_re_out(1563),
            product_im_out=>mul_im_out(1563)
        );

    UMUL_1564 : complex_multiplier
    generic map(
            re_multiplicator=>-9102, --- -0.555541992188 + j0.831420898438
            im_multiplicator=>13622
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1564),
            data_im_in=>first_stage_im_out(1564),
            product_re_out=>mul_re_out(1564),
            product_im_out=>mul_im_out(1564)
        );

    UMUL_1565 : complex_multiplier
    generic map(
            re_multiplicator=>-7005, --- -0.427551269531 + j0.903930664062
            im_multiplicator=>14810
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1565),
            data_im_in=>first_stage_im_out(1565),
            product_re_out=>mul_re_out(1565),
            product_im_out=>mul_im_out(1565)
        );

    UMUL_1566 : complex_multiplier
    generic map(
            re_multiplicator=>-4756, --- -0.290283203125 + j0.956909179688
            im_multiplicator=>15678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1566),
            data_im_in=>first_stage_im_out(1566),
            product_re_out=>mul_re_out(1566),
            product_im_out=>mul_im_out(1566)
        );

    UMUL_1567 : complex_multiplier
    generic map(
            re_multiplicator=>-2404, --- -0.146728515625 + j0.989135742188
            im_multiplicator=>16206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1567),
            data_im_in=>first_stage_im_out(1567),
            product_re_out=>mul_re_out(1567),
            product_im_out=>mul_im_out(1567)
        );

    UDELAY_1568_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1568),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1568)
        );
    UDELAY_1568_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1568),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1568)
        );
    USHIFTER_1568_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1568),
            data_out=>mul_re_out(1568)
        );
    USHIFTER_1568_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1568),
            data_out=>mul_im_out(1568)
        );

    UMUL_1569 : complex_multiplier
    generic map(
            re_multiplicator=>16199, --- 0.988708496094 + j-0.149719238281
            im_multiplicator=>-2453
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1569),
            data_im_in=>first_stage_im_out(1569),
            product_re_out=>mul_re_out(1569),
            product_im_out=>mul_im_out(1569)
        );

    UMUL_1570 : complex_multiplier
    generic map(
            re_multiplicator=>15649, --- 0.955139160156 + j-0.296142578125
            im_multiplicator=>-4852
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1570),
            data_im_in=>first_stage_im_out(1570),
            product_re_out=>mul_re_out(1570),
            product_im_out=>mul_im_out(1570)
        );

    UMUL_1571 : complex_multiplier
    generic map(
            re_multiplicator=>14745, --- 0.899963378906 + j-0.435852050781
            im_multiplicator=>-7141
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1571),
            data_im_in=>first_stage_im_out(1571),
            product_re_out=>mul_re_out(1571),
            product_im_out=>mul_im_out(1571)
        );

    UMUL_1572 : complex_multiplier
    generic map(
            re_multiplicator=>13510, --- 0.824584960938 + j-0.565673828125
            im_multiplicator=>-9268
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1572),
            data_im_in=>first_stage_im_out(1572),
            product_re_out=>mul_re_out(1572),
            product_im_out=>mul_im_out(1572)
        );

    UMUL_1573 : complex_multiplier
    generic map(
            re_multiplicator=>11969, --- 0.730529785156 + j-0.682800292969
            im_multiplicator=>-11187
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1573),
            data_im_in=>first_stage_im_out(1573),
            product_re_out=>mul_re_out(1573),
            product_im_out=>mul_im_out(1573)
        );

    UMUL_1574 : complex_multiplier
    generic map(
            re_multiplicator=>10159, --- 0.620056152344 + j-0.784545898438
            im_multiplicator=>-12854
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1574),
            data_im_in=>first_stage_im_out(1574),
            product_re_out=>mul_re_out(1574),
            product_im_out=>mul_im_out(1574)
        );

    UMUL_1575 : complex_multiplier
    generic map(
            re_multiplicator=>8119, --- 0.495544433594 + j-0.868530273438
            im_multiplicator=>-14230
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1575),
            data_im_in=>first_stage_im_out(1575),
            product_re_out=>mul_re_out(1575),
            product_im_out=>mul_im_out(1575)
        );

    UMUL_1576 : complex_multiplier
    generic map(
            re_multiplicator=>5896, --- 0.35986328125 + j-0.932983398438
            im_multiplicator=>-15286
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1576),
            data_im_in=>first_stage_im_out(1576),
            product_re_out=>mul_re_out(1576),
            product_im_out=>mul_im_out(1576)
        );

    UMUL_1577 : complex_multiplier
    generic map(
            re_multiplicator=>3540, --- 0.216064453125 + j-0.976318359375
            im_multiplicator=>-15996
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1577),
            data_im_in=>first_stage_im_out(1577),
            product_re_out=>mul_re_out(1577),
            product_im_out=>mul_im_out(1577)
        );

    UMUL_1578 : complex_multiplier
    generic map(
            re_multiplicator=>1105, --- 0.0674438476562 + j-0.997680664062
            im_multiplicator=>-16346
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1578),
            data_im_in=>first_stage_im_out(1578),
            product_re_out=>mul_re_out(1578),
            product_im_out=>mul_im_out(1578)
        );

    UMUL_1579 : complex_multiplier
    generic map(
            re_multiplicator=>-1355, --- -0.0827026367188 + j-0.996520996094
            im_multiplicator=>-16327
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1579),
            data_im_in=>first_stage_im_out(1579),
            product_re_out=>mul_re_out(1579),
            product_im_out=>mul_im_out(1579)
        );

    UMUL_1580 : complex_multiplier
    generic map(
            re_multiplicator=>-3785, --- -0.231018066406 + j-0.972900390625
            im_multiplicator=>-15940
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1580),
            data_im_in=>first_stage_im_out(1580),
            product_re_out=>mul_re_out(1580),
            product_im_out=>mul_im_out(1580)
        );

    UMUL_1581 : complex_multiplier
    generic map(
            re_multiplicator=>-6130, --- -0.374145507812 + j-0.927307128906
            im_multiplicator=>-15193
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1581),
            data_im_in=>first_stage_im_out(1581),
            product_re_out=>mul_re_out(1581),
            product_im_out=>mul_im_out(1581)
        );

    UMUL_1582 : complex_multiplier
    generic map(
            re_multiplicator=>-8336, --- -0.5087890625 + j-0.86083984375
            im_multiplicator=>-14104
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1582),
            data_im_in=>first_stage_im_out(1582),
            product_re_out=>mul_re_out(1582),
            product_im_out=>mul_im_out(1582)
        );

    UMUL_1583 : complex_multiplier
    generic map(
            re_multiplicator=>-10354, --- -0.631958007812 + j-0.77490234375
            im_multiplicator=>-12696
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1583),
            data_im_in=>first_stage_im_out(1583),
            product_re_out=>mul_re_out(1583),
            product_im_out=>mul_im_out(1583)
        );

    UMUL_1584 : complex_multiplier
    generic map(
            re_multiplicator=>-12139, --- -0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1584),
            data_im_in=>first_stage_im_out(1584),
            product_re_out=>mul_re_out(1584),
            product_im_out=>mul_im_out(1584)
        );

    UMUL_1585 : complex_multiplier
    generic map(
            re_multiplicator=>-13650, --- -0.833129882812 + j-0.552978515625
            im_multiplicator=>-9060
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1585),
            data_im_in=>first_stage_im_out(1585),
            product_re_out=>mul_re_out(1585),
            product_im_out=>mul_im_out(1585)
        );

    UMUL_1586 : complex_multiplier
    generic map(
            re_multiplicator=>-14853, --- -0.906555175781 + j-0.421997070312
            im_multiplicator=>-6914
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1586),
            data_im_in=>first_stage_im_out(1586),
            product_re_out=>mul_re_out(1586),
            product_im_out=>mul_im_out(1586)
        );

    UMUL_1587 : complex_multiplier
    generic map(
            re_multiplicator=>-15721, --- -0.959533691406 + j-0.281433105469
            im_multiplicator=>-4611
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1587),
            data_im_in=>first_stage_im_out(1587),
            product_re_out=>mul_re_out(1587),
            product_im_out=>mul_im_out(1587)
        );

    UMUL_1588 : complex_multiplier
    generic map(
            re_multiplicator=>-16234, --- -0.990844726562 + j-0.134521484375
            im_multiplicator=>-2204
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1588),
            data_im_in=>first_stage_im_out(1588),
            product_re_out=>mul_re_out(1588),
            product_im_out=>mul_im_out(1588)
        );

    UMUL_1589 : complex_multiplier
    generic map(
            re_multiplicator=>-16382, --- -0.999877929688 + j0.0153198242188
            im_multiplicator=>251
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1589),
            data_im_in=>first_stage_im_out(1589),
            product_re_out=>mul_re_out(1589),
            product_im_out=>mul_im_out(1589)
        );

    UMUL_1590 : complex_multiplier
    generic map(
            re_multiplicator=>-16159, --- -0.986267089844 + j0.164855957031
            im_multiplicator=>2701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1590),
            data_im_in=>first_stage_im_out(1590),
            product_re_out=>mul_re_out(1590),
            product_im_out=>mul_im_out(1590)
        );

    UMUL_1591 : complex_multiplier
    generic map(
            re_multiplicator=>-15572, --- -0.950439453125 + j0.310729980469
            im_multiplicator=>5091
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1591),
            data_im_in=>first_stage_im_out(1591),
            product_re_out=>mul_re_out(1591),
            product_im_out=>mul_im_out(1591)
        );

    UMUL_1592 : complex_multiplier
    generic map(
            re_multiplicator=>-14634, --- -0.893188476562 + j0.449584960938
            im_multiplicator=>7366
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1592),
            data_im_in=>first_stage_im_out(1592),
            product_re_out=>mul_re_out(1592),
            product_im_out=>mul_im_out(1592)
        );

    UMUL_1593 : complex_multiplier
    generic map(
            re_multiplicator=>-13366, --- -0.815795898438 + j0.578308105469
            im_multiplicator=>9475
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1593),
            data_im_in=>first_stage_im_out(1593),
            product_re_out=>mul_re_out(1593),
            product_im_out=>mul_im_out(1593)
        );

    UMUL_1594 : complex_multiplier
    generic map(
            re_multiplicator=>-11796, --- -0.719970703125 + j0.693969726562
            im_multiplicator=>11370
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1594),
            data_im_in=>first_stage_im_out(1594),
            product_re_out=>mul_re_out(1594),
            product_im_out=>mul_im_out(1594)
        );

    UMUL_1595 : complex_multiplier
    generic map(
            re_multiplicator=>-9960, --- -0.60791015625 + j0.7939453125
            im_multiplicator=>13008
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1595),
            data_im_in=>first_stage_im_out(1595),
            product_re_out=>mul_re_out(1595),
            product_im_out=>mul_im_out(1595)
        );

    UMUL_1596 : complex_multiplier
    generic map(
            re_multiplicator=>-7900, --- -0.482177734375 + j0.876037597656
            im_multiplicator=>14353
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1596),
            data_im_in=>first_stage_im_out(1596),
            product_re_out=>mul_re_out(1596),
            product_im_out=>mul_im_out(1596)
        );

    UMUL_1597 : complex_multiplier
    generic map(
            re_multiplicator=>-5661, --- -0.345520019531 + j0.938354492188
            im_multiplicator=>15374
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1597),
            data_im_in=>first_stage_im_out(1597),
            product_re_out=>mul_re_out(1597),
            product_im_out=>mul_im_out(1597)
        );

    UMUL_1598 : complex_multiplier
    generic map(
            re_multiplicator=>-3294, --- -0.201049804688 + j0.979553222656
            im_multiplicator=>16049
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1598),
            data_im_in=>first_stage_im_out(1598),
            product_re_out=>mul_re_out(1598),
            product_im_out=>mul_im_out(1598)
        );

    UMUL_1599 : complex_multiplier
    generic map(
            re_multiplicator=>-854, --- -0.0521240234375 + j0.998596191406
            im_multiplicator=>16361
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1599),
            data_im_in=>first_stage_im_out(1599),
            product_re_out=>mul_re_out(1599),
            product_im_out=>mul_im_out(1599)
        );

    UDELAY_1600_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1600),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1600)
        );
    UDELAY_1600_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1600),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1600)
        );
    USHIFTER_1600_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1600),
            data_out=>mul_re_out(1600)
        );
    USHIFTER_1600_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1600),
            data_out=>mul_im_out(1600)
        );

    UMUL_1601 : complex_multiplier
    generic map(
            re_multiplicator=>16191, --- 0.988220214844 + j-0.152770996094
            im_multiplicator=>-2503
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1601),
            data_im_in=>first_stage_im_out(1601),
            product_re_out=>mul_re_out(1601),
            product_im_out=>mul_im_out(1601)
        );

    UMUL_1602 : complex_multiplier
    generic map(
            re_multiplicator=>15618, --- 0.953247070312 + j-0.302001953125
            im_multiplicator=>-4948
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1602),
            data_im_in=>first_stage_im_out(1602),
            product_re_out=>mul_re_out(1602),
            product_im_out=>mul_im_out(1602)
        );

    UMUL_1603 : complex_multiplier
    generic map(
            re_multiplicator=>14679, --- 0.895935058594 + j-0.444091796875
            im_multiplicator=>-7276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1603),
            data_im_in=>first_stage_im_out(1603),
            product_re_out=>mul_re_out(1603),
            product_im_out=>mul_im_out(1603)
        );

    UMUL_1604 : complex_multiplier
    generic map(
            re_multiplicator=>13395, --- 0.817565917969 + j-0.575805664062
            im_multiplicator=>-9434
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1604),
            data_im_in=>first_stage_im_out(1604),
            product_re_out=>mul_re_out(1604),
            product_im_out=>mul_im_out(1604)
        );

    UMUL_1605 : complex_multiplier
    generic map(
            re_multiplicator=>11796, --- 0.719970703125 + j-0.693969726562
            im_multiplicator=>-11370
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1605),
            data_im_in=>first_stage_im_out(1605),
            product_re_out=>mul_re_out(1605),
            product_im_out=>mul_im_out(1605)
        );

    UMUL_1606 : complex_multiplier
    generic map(
            re_multiplicator=>9920, --- 0.60546875 + j-0.795776367188
            im_multiplicator=>-13038
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1606),
            data_im_in=>first_stage_im_out(1606),
            product_re_out=>mul_re_out(1606),
            product_im_out=>mul_im_out(1606)
        );

    UMUL_1607 : complex_multiplier
    generic map(
            re_multiplicator=>7811, --- 0.476745605469 + j-0.878967285156
            im_multiplicator=>-14401
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1607),
            data_im_in=>first_stage_im_out(1607),
            product_re_out=>mul_re_out(1607),
            product_im_out=>mul_im_out(1607)
        );

    UMUL_1608 : complex_multiplier
    generic map(
            re_multiplicator=>5519, --- 0.336853027344 + j-0.941528320312
            im_multiplicator=>-15426
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1608),
            data_im_in=>first_stage_im_out(1608),
            product_re_out=>mul_re_out(1608),
            product_im_out=>mul_im_out(1608)
        );

    UMUL_1609 : complex_multiplier
    generic map(
            re_multiplicator=>3097, --- 0.189025878906 + j-0.98193359375
            im_multiplicator=>-16088
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1609),
            data_im_in=>first_stage_im_out(1609),
            product_re_out=>mul_re_out(1609),
            product_im_out=>mul_im_out(1609)
        );

    UMUL_1610 : complex_multiplier
    generic map(
            re_multiplicator=>603, --- 0.0368041992188 + j-0.999267578125
            im_multiplicator=>-16372
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1610),
            data_im_in=>first_stage_im_out(1610),
            product_re_out=>mul_re_out(1610),
            product_im_out=>mul_im_out(1610)
        );

    UMUL_1611 : complex_multiplier
    generic map(
            re_multiplicator=>-1905, --- -0.116271972656 + j-0.9931640625
            im_multiplicator=>-16272
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1611),
            data_im_in=>first_stage_im_out(1611),
            product_re_out=>mul_re_out(1611),
            product_im_out=>mul_im_out(1611)
        );

    UMUL_1612 : complex_multiplier
    generic map(
            re_multiplicator=>-4369, --- -0.266662597656 + j-0.963745117188
            im_multiplicator=>-15790
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1612),
            data_im_in=>first_stage_im_out(1612),
            product_re_out=>mul_re_out(1612),
            product_im_out=>mul_im_out(1612)
        );

    UMUL_1613 : complex_multiplier
    generic map(
            re_multiplicator=>-6731, --- -0.410827636719 + j-0.911682128906
            im_multiplicator=>-14937
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1613),
            data_im_in=>first_stage_im_out(1613),
            product_re_out=>mul_re_out(1613),
            product_im_out=>mul_im_out(1613)
        );

    UMUL_1614 : complex_multiplier
    generic map(
            re_multiplicator=>-8934, --- -0.545288085938 + j-0.838195800781
            im_multiplicator=>-13733
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1614),
            data_im_in=>first_stage_im_out(1614),
            product_re_out=>mul_re_out(1614),
            product_im_out=>mul_im_out(1614)
        );

    UMUL_1615 : complex_multiplier
    generic map(
            re_multiplicator=>-10928, --- -0.6669921875 + j-0.745056152344
            im_multiplicator=>-12207
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1615),
            data_im_in=>first_stage_im_out(1615),
            product_re_out=>mul_re_out(1615),
            product_im_out=>mul_im_out(1615)
        );

    UMUL_1616 : complex_multiplier
    generic map(
            re_multiplicator=>-12665, --- -0.773010253906 + j-0.634338378906
            im_multiplicator=>-10393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1616),
            data_im_in=>first_stage_im_out(1616),
            product_re_out=>mul_re_out(1616),
            product_im_out=>mul_im_out(1616)
        );

    UMUL_1617 : complex_multiplier
    generic map(
            re_multiplicator=>-14104, --- -0.86083984375 + j-0.5087890625
            im_multiplicator=>-8336
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1617),
            data_im_in=>first_stage_im_out(1617),
            product_re_out=>mul_re_out(1617),
            product_im_out=>mul_im_out(1617)
        );

    UMUL_1618 : complex_multiplier
    generic map(
            re_multiplicator=>-15212, --- -0.928466796875 + j-0.371276855469
            im_multiplicator=>-6083
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1618),
            data_im_in=>first_stage_im_out(1618),
            product_re_out=>mul_re_out(1618),
            product_im_out=>mul_im_out(1618)
        );

    UMUL_1619 : complex_multiplier
    generic map(
            re_multiplicator=>-15963, --- -0.974304199219 + j-0.225036621094
            im_multiplicator=>-3687
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1619),
            data_im_in=>first_stage_im_out(1619),
            product_re_out=>mul_re_out(1619),
            product_im_out=>mul_im_out(1619)
        );

    UMUL_1620 : complex_multiplier
    generic map(
            re_multiplicator=>-16339, --- -0.997253417969 + j-0.0735473632812
            im_multiplicator=>-1205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1620),
            data_im_in=>first_stage_im_out(1620),
            product_re_out=>mul_re_out(1620),
            product_im_out=>mul_im_out(1620)
        );

    UMUL_1621 : complex_multiplier
    generic map(
            re_multiplicator=>-16331, --- -0.996765136719 + j0.0796508789062
            im_multiplicator=>1305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1621),
            data_im_in=>first_stage_im_out(1621),
            product_re_out=>mul_re_out(1621),
            product_im_out=>mul_im_out(1621)
        );

    UMUL_1622 : complex_multiplier
    generic map(
            re_multiplicator=>-15940, --- -0.972900390625 + j0.231018066406
            im_multiplicator=>3785
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1622),
            data_im_in=>first_stage_im_out(1622),
            product_re_out=>mul_re_out(1622),
            product_im_out=>mul_im_out(1622)
        );

    UMUL_1623 : complex_multiplier
    generic map(
            re_multiplicator=>-15175, --- -0.926208496094 + j0.376953125
            im_multiplicator=>6176
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1623),
            data_im_in=>first_stage_im_out(1623),
            product_re_out=>mul_re_out(1623),
            product_im_out=>mul_im_out(1623)
        );

    UMUL_1624 : complex_multiplier
    generic map(
            re_multiplicator=>-14053, --- -0.857727050781 + j0.514099121094
            im_multiplicator=>8423
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1624),
            data_im_in=>first_stage_im_out(1624),
            product_re_out=>mul_re_out(1624),
            product_im_out=>mul_im_out(1624)
        );

    UMUL_1625 : complex_multiplier
    generic map(
            re_multiplicator=>-12600, --- -0.76904296875 + j0.639099121094
            im_multiplicator=>10471
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1625),
            data_im_in=>first_stage_im_out(1625),
            product_re_out=>mul_re_out(1625),
            product_im_out=>mul_im_out(1625)
        );

    UMUL_1626 : complex_multiplier
    generic map(
            re_multiplicator=>-10853, --- -0.662414550781 + j0.749084472656
            im_multiplicator=>12273
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1626),
            data_im_in=>first_stage_im_out(1626),
            product_re_out=>mul_re_out(1626),
            product_im_out=>mul_im_out(1626)
        );

    UMUL_1627 : complex_multiplier
    generic map(
            re_multiplicator=>-8850, --- -0.540161132812 + j0.841552734375
            im_multiplicator=>13788
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1627),
            data_im_in=>first_stage_im_out(1627),
            product_re_out=>mul_re_out(1627),
            product_im_out=>mul_im_out(1627)
        );

    UMUL_1628 : complex_multiplier
    generic map(
            re_multiplicator=>-6639, --- -0.405212402344 + j0.914184570312
            im_multiplicator=>14978
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1628),
            data_im_in=>first_stage_im_out(1628),
            product_re_out=>mul_re_out(1628),
            product_im_out=>mul_im_out(1628)
        );

    UMUL_1629 : complex_multiplier
    generic map(
            re_multiplicator=>-4272, --- -0.2607421875 + j0.965393066406
            im_multiplicator=>15817
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1629),
            data_im_in=>first_stage_im_out(1629),
            product_re_out=>mul_re_out(1629),
            product_im_out=>mul_im_out(1629)
        );

    UMUL_1630 : complex_multiplier
    generic map(
            re_multiplicator=>-1805, --- -0.110168457031 + j0.993896484375
            im_multiplicator=>16284
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1630),
            data_im_in=>first_stage_im_out(1630),
            product_re_out=>mul_re_out(1630),
            product_im_out=>mul_im_out(1630)
        );

    UMUL_1631 : complex_multiplier
    generic map(
            re_multiplicator=>703, --- 0.0429077148438 + j0.9990234375
            im_multiplicator=>16368
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1631),
            data_im_in=>first_stage_im_out(1631),
            product_re_out=>mul_re_out(1631),
            product_im_out=>mul_im_out(1631)
        );

    UDELAY_1632_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1632),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1632)
        );
    UDELAY_1632_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1632),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1632)
        );
    USHIFTER_1632_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1632),
            data_out=>mul_re_out(1632)
        );
    USHIFTER_1632_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1632),
            data_out=>mul_im_out(1632)
        );

    UMUL_1633 : complex_multiplier
    generic map(
            re_multiplicator=>16183, --- 0.987731933594 + j-0.155822753906
            im_multiplicator=>-2553
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1633),
            data_im_in=>first_stage_im_out(1633),
            product_re_out=>mul_re_out(1633),
            product_im_out=>mul_im_out(1633)
        );

    UMUL_1634 : complex_multiplier
    generic map(
            re_multiplicator=>15588, --- 0.951416015625 + j-0.307800292969
            im_multiplicator=>-5043
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1634),
            data_im_in=>first_stage_im_out(1634),
            product_re_out=>mul_re_out(1634),
            product_im_out=>mul_im_out(1634)
        );

    UMUL_1635 : complex_multiplier
    generic map(
            re_multiplicator=>14611, --- 0.891784667969 + j-0.452331542969
            im_multiplicator=>-7411
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1635),
            data_im_in=>first_stage_im_out(1635),
            product_re_out=>mul_re_out(1635),
            product_im_out=>mul_im_out(1635)
        );

    UMUL_1636 : complex_multiplier
    generic map(
            re_multiplicator=>13278, --- 0.810424804688 + j-0.585754394531
            im_multiplicator=>-9597
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1636),
            data_im_in=>first_stage_im_out(1636),
            product_re_out=>mul_re_out(1636),
            product_im_out=>mul_im_out(1636)
        );

    UMUL_1637 : complex_multiplier
    generic map(
            re_multiplicator=>11620, --- 0.709228515625 + j-0.704895019531
            im_multiplicator=>-11549
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1637),
            data_im_in=>first_stage_im_out(1637),
            product_re_out=>mul_re_out(1637),
            product_im_out=>mul_im_out(1637)
        );

    UMUL_1638 : complex_multiplier
    generic map(
            re_multiplicator=>9679, --- 0.590759277344 + j-0.806823730469
            im_multiplicator=>-13219
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1638),
            data_im_in=>first_stage_im_out(1638),
            product_re_out=>mul_re_out(1638),
            product_im_out=>mul_im_out(1638)
        );

    UMUL_1639 : complex_multiplier
    generic map(
            re_multiplicator=>7500, --- 0.457763671875 + j-0.889038085938
            im_multiplicator=>-14566
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1639),
            data_im_in=>first_stage_im_out(1639),
            product_re_out=>mul_re_out(1639),
            product_im_out=>mul_im_out(1639)
        );

    UMUL_1640 : complex_multiplier
    generic map(
            re_multiplicator=>5139, --- 0.313659667969 + j-0.949523925781
            im_multiplicator=>-15557
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1640),
            data_im_in=>first_stage_im_out(1640),
            product_re_out=>mul_re_out(1640),
            product_im_out=>mul_im_out(1640)
        );

    UMUL_1641 : complex_multiplier
    generic map(
            re_multiplicator=>2652, --- 0.161865234375 + j-0.986755371094
            im_multiplicator=>-16167
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1641),
            data_im_in=>first_stage_im_out(1641),
            product_re_out=>mul_re_out(1641),
            product_im_out=>mul_im_out(1641)
        );

    UMUL_1642 : complex_multiplier
    generic map(
            re_multiplicator=>100, --- 0.006103515625 + j-0.999938964844
            im_multiplicator=>-16383
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1642),
            data_im_in=>first_stage_im_out(1642),
            product_re_out=>mul_re_out(1642),
            product_im_out=>mul_im_out(1642)
        );

    UMUL_1643 : complex_multiplier
    generic map(
            re_multiplicator=>-2453, --- -0.149719238281 + j-0.988708496094
            im_multiplicator=>-16199
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1643),
            data_im_in=>first_stage_im_out(1643),
            product_re_out=>mul_re_out(1643),
            product_im_out=>mul_im_out(1643)
        );

    UMUL_1644 : complex_multiplier
    generic map(
            re_multiplicator=>-4948, --- -0.302001953125 + j-0.953247070312
            im_multiplicator=>-15618
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1644),
            data_im_in=>first_stage_im_out(1644),
            product_re_out=>mul_re_out(1644),
            product_im_out=>mul_im_out(1644)
        );

    UMUL_1645 : complex_multiplier
    generic map(
            re_multiplicator=>-7321, --- -0.446838378906 + j-0.894592285156
            im_multiplicator=>-14657
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1645),
            data_im_in=>first_stage_im_out(1645),
            product_re_out=>mul_re_out(1645),
            product_im_out=>mul_im_out(1645)
        );

    UMUL_1646 : complex_multiplier
    generic map(
            re_multiplicator=>-9516, --- -0.580810546875 + j-0.814025878906
            im_multiplicator=>-13337
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1646),
            data_im_in=>first_stage_im_out(1646),
            product_re_out=>mul_re_out(1646),
            product_im_out=>mul_im_out(1646)
        );

    UMUL_1647 : complex_multiplier
    generic map(
            re_multiplicator=>-11478, --- -0.700561523438 + j-0.713562011719
            im_multiplicator=>-11691
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1647),
            data_im_in=>first_stage_im_out(1647),
            product_re_out=>mul_re_out(1647),
            product_im_out=>mul_im_out(1647)
        );

    UMUL_1648 : complex_multiplier
    generic map(
            re_multiplicator=>-13159, --- -0.803161621094 + j-0.595642089844
            im_multiplicator=>-9759
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1648),
            data_im_in=>first_stage_im_out(1648),
            product_re_out=>mul_re_out(1648),
            product_im_out=>mul_im_out(1648)
        );

    UMUL_1649 : complex_multiplier
    generic map(
            re_multiplicator=>-14519, --- -0.886169433594 + j-0.463256835938
            im_multiplicator=>-7590
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1649),
            data_im_in=>first_stage_im_out(1649),
            product_re_out=>mul_re_out(1649),
            product_im_out=>mul_im_out(1649)
        );

    UMUL_1650 : complex_multiplier
    generic map(
            re_multiplicator=>-15525, --- -0.947570800781 + j-0.319458007812
            im_multiplicator=>-5234
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1650),
            data_im_in=>first_stage_im_out(1650),
            product_re_out=>mul_re_out(1650),
            product_im_out=>mul_im_out(1650)
        );

    UMUL_1651 : complex_multiplier
    generic map(
            re_multiplicator=>-16151, --- -0.985778808594 + j-0.167907714844
            im_multiplicator=>-2751
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1651),
            data_im_in=>first_stage_im_out(1651),
            product_re_out=>mul_re_out(1651),
            product_im_out=>mul_im_out(1651)
        );

    UMUL_1652 : complex_multiplier
    generic map(
            re_multiplicator=>-16382, --- -0.999877929688 + j-0.0122680664062
            im_multiplicator=>-201
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1652),
            data_im_in=>first_stage_im_out(1652),
            product_re_out=>mul_re_out(1652),
            product_im_out=>mul_im_out(1652)
        );

    UMUL_1653 : complex_multiplier
    generic map(
            re_multiplicator=>-16213, --- -0.989562988281 + j0.143676757812
            im_multiplicator=>2354
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1653),
            data_im_in=>first_stage_im_out(1653),
            product_re_out=>mul_re_out(1653),
            product_im_out=>mul_im_out(1653)
        );

    UMUL_1654 : complex_multiplier
    generic map(
            re_multiplicator=>-15649, --- -0.955139160156 + j0.296142578125
            im_multiplicator=>4852
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1654),
            data_im_in=>first_stage_im_out(1654),
            product_re_out=>mul_re_out(1654),
            product_im_out=>mul_im_out(1654)
        );

    UMUL_1655 : complex_multiplier
    generic map(
            re_multiplicator=>-14701, --- -0.897277832031 + j0.441345214844
            im_multiplicator=>7231
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1655),
            data_im_in=>first_stage_im_out(1655),
            product_re_out=>mul_re_out(1655),
            product_im_out=>mul_im_out(1655)
        );

    UMUL_1656 : complex_multiplier
    generic map(
            re_multiplicator=>-13395, --- -0.817565917969 + j0.575805664062
            im_multiplicator=>9434
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1656),
            data_im_in=>first_stage_im_out(1656),
            product_re_out=>mul_re_out(1656),
            product_im_out=>mul_im_out(1656)
        );

    UMUL_1657 : complex_multiplier
    generic map(
            re_multiplicator=>-11761, --- -0.717834472656 + j0.696166992188
            im_multiplicator=>11406
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1657),
            data_im_in=>first_stage_im_out(1657),
            product_re_out=>mul_re_out(1657),
            product_im_out=>mul_im_out(1657)
        );

    UMUL_1658 : complex_multiplier
    generic map(
            re_multiplicator=>-9840, --- -0.6005859375 + j0.799499511719
            im_multiplicator=>13099
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1658),
            data_im_in=>first_stage_im_out(1658),
            product_re_out=>mul_re_out(1658),
            product_im_out=>mul_im_out(1658)
        );

    UMUL_1659 : complex_multiplier
    generic map(
            re_multiplicator=>-7678, --- -0.468627929688 + j0.883361816406
            im_multiplicator=>14473
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1659),
            data_im_in=>first_stage_im_out(1659),
            product_re_out=>mul_re_out(1659),
            product_im_out=>mul_im_out(1659)
        );

    UMUL_1660 : complex_multiplier
    generic map(
            re_multiplicator=>-5329, --- -0.325256347656 + j0.945556640625
            im_multiplicator=>15492
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1660),
            data_im_in=>first_stage_im_out(1660),
            product_re_out=>mul_re_out(1660),
            product_im_out=>mul_im_out(1660)
        );

    UMUL_1661 : complex_multiplier
    generic map(
            re_multiplicator=>-2850, --- -0.173950195312 + j0.984741210938
            im_multiplicator=>16134
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1661),
            data_im_in=>first_stage_im_out(1661),
            product_re_out=>mul_re_out(1661),
            product_im_out=>mul_im_out(1661)
        );

    UMUL_1662 : complex_multiplier
    generic map(
            re_multiplicator=>-301, --- -0.0183715820312 + j0.999816894531
            im_multiplicator=>16381
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1662),
            data_im_in=>first_stage_im_out(1662),
            product_re_out=>mul_re_out(1662),
            product_im_out=>mul_im_out(1662)
        );

    UMUL_1663 : complex_multiplier
    generic map(
            re_multiplicator=>2254, --- 0.137573242188 + j0.990478515625
            im_multiplicator=>16228
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1663),
            data_im_in=>first_stage_im_out(1663),
            product_re_out=>mul_re_out(1663),
            product_im_out=>mul_im_out(1663)
        );

    UDELAY_1664_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1664),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1664)
        );
    UDELAY_1664_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1664),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1664)
        );
    USHIFTER_1664_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1664),
            data_out=>mul_re_out(1664)
        );
    USHIFTER_1664_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1664),
            data_out=>mul_im_out(1664)
        );

    UMUL_1665 : complex_multiplier
    generic map(
            re_multiplicator=>16175, --- 0.987243652344 + j-0.158813476562
            im_multiplicator=>-2602
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1665),
            data_im_in=>first_stage_im_out(1665),
            product_re_out=>mul_re_out(1665),
            product_im_out=>mul_im_out(1665)
        );

    UMUL_1666 : complex_multiplier
    generic map(
            re_multiplicator=>15557, --- 0.949523925781 + j-0.313659667969
            im_multiplicator=>-5139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1666),
            data_im_in=>first_stage_im_out(1666),
            product_re_out=>mul_re_out(1666),
            product_im_out=>mul_im_out(1666)
        );

    UMUL_1667 : complex_multiplier
    generic map(
            re_multiplicator=>14543, --- 0.887634277344 + j-0.460510253906
            im_multiplicator=>-7545
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1667),
            data_im_in=>first_stage_im_out(1667),
            product_re_out=>mul_re_out(1667),
            product_im_out=>mul_im_out(1667)
        );

    UMUL_1668 : complex_multiplier
    generic map(
            re_multiplicator=>13159, --- 0.803161621094 + j-0.595642089844
            im_multiplicator=>-9759
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1668),
            data_im_in=>first_stage_im_out(1668),
            product_re_out=>mul_re_out(1668),
            product_im_out=>mul_im_out(1668)
        );

    UMUL_1669 : complex_multiplier
    generic map(
            re_multiplicator=>11442, --- 0.698364257812 + j-0.715698242188
            im_multiplicator=>-11726
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1669),
            data_im_in=>first_stage_im_out(1669),
            product_re_out=>mul_re_out(1669),
            product_im_out=>mul_im_out(1669)
        );

    UMUL_1670 : complex_multiplier
    generic map(
            re_multiplicator=>9434, --- 0.575805664062 + j-0.817565917969
            im_multiplicator=>-13395
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1670),
            data_im_in=>first_stage_im_out(1670),
            product_re_out=>mul_re_out(1670),
            product_im_out=>mul_im_out(1670)
        );

    UMUL_1671 : complex_multiplier
    generic map(
            re_multiplicator=>7186, --- 0.438598632812 + j-0.898620605469
            im_multiplicator=>-14723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1671),
            data_im_in=>first_stage_im_out(1671),
            product_re_out=>mul_re_out(1671),
            product_im_out=>mul_im_out(1671)
        );

    UMUL_1672 : complex_multiplier
    generic map(
            re_multiplicator=>4756, --- 0.290283203125 + j-0.956909179688
            im_multiplicator=>-15678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1672),
            data_im_in=>first_stage_im_out(1672),
            product_re_out=>mul_re_out(1672),
            product_im_out=>mul_im_out(1672)
        );

    UMUL_1673 : complex_multiplier
    generic map(
            re_multiplicator=>2204, --- 0.134521484375 + j-0.990844726562
            im_multiplicator=>-16234
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1673),
            data_im_in=>first_stage_im_out(1673),
            product_re_out=>mul_re_out(1673),
            product_im_out=>mul_im_out(1673)
        );

    UMUL_1674 : complex_multiplier
    generic map(
            re_multiplicator=>-402, --- -0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1674),
            data_im_in=>first_stage_im_out(1674),
            product_re_out=>mul_re_out(1674),
            product_im_out=>mul_im_out(1674)
        );

    UMUL_1675 : complex_multiplier
    generic map(
            re_multiplicator=>-2998, --- -0.182983398438 + j-0.983093261719
            im_multiplicator=>-16107
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1675),
            data_im_in=>first_stage_im_out(1675),
            product_re_out=>mul_re_out(1675),
            product_im_out=>mul_im_out(1675)
        );

    UMUL_1676 : complex_multiplier
    generic map(
            re_multiplicator=>-5519, --- -0.336853027344 + j-0.941528320312
            im_multiplicator=>-15426
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1676),
            data_im_in=>first_stage_im_out(1676),
            product_re_out=>mul_re_out(1676),
            product_im_out=>mul_im_out(1676)
        );

    UMUL_1677 : complex_multiplier
    generic map(
            re_multiplicator=>-7900, --- -0.482177734375 + j-0.876037597656
            im_multiplicator=>-14353
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1677),
            data_im_in=>first_stage_im_out(1677),
            product_re_out=>mul_re_out(1677),
            product_im_out=>mul_im_out(1677)
        );

    UMUL_1678 : complex_multiplier
    generic map(
            re_multiplicator=>-10079, --- -0.615173339844 + j-0.788330078125
            im_multiplicator=>-12916
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1678),
            data_im_in=>first_stage_im_out(1678),
            product_re_out=>mul_re_out(1678),
            product_im_out=>mul_im_out(1678)
        );

    UMUL_1679 : complex_multiplier
    generic map(
            re_multiplicator=>-12003, --- -0.732604980469 + j-0.680541992188
            im_multiplicator=>-11150
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1679),
            data_im_in=>first_stage_im_out(1679),
            product_re_out=>mul_re_out(1679),
            product_im_out=>mul_im_out(1679)
        );

    UMUL_1680 : complex_multiplier
    generic map(
            re_multiplicator=>-13622, --- -0.831420898438 + j-0.555541992188
            im_multiplicator=>-9102
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1680),
            data_im_in=>first_stage_im_out(1680),
            product_re_out=>mul_re_out(1680),
            product_im_out=>mul_im_out(1680)
        );

    UMUL_1681 : complex_multiplier
    generic map(
            re_multiplicator=>-14895, --- -0.909118652344 + j-0.416381835938
            im_multiplicator=>-6822
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1681),
            data_im_in=>first_stage_im_out(1681),
            product_re_out=>mul_re_out(1681),
            product_im_out=>mul_im_out(1681)
        );

    UMUL_1682 : complex_multiplier
    generic map(
            re_multiplicator=>-15790, --- -0.963745117188 + j-0.266662597656
            im_multiplicator=>-4369
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1682),
            data_im_in=>first_stage_im_out(1682),
            product_re_out=>mul_re_out(1682),
            product_im_out=>mul_im_out(1682)
        );

    UMUL_1683 : complex_multiplier
    generic map(
            re_multiplicator=>-16284, --- -0.993896484375 + j-0.110168457031
            im_multiplicator=>-1805
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1683),
            data_im_in=>first_stage_im_out(1683),
            product_re_out=>mul_re_out(1683),
            product_im_out=>mul_im_out(1683)
        );

    UMUL_1684 : complex_multiplier
    generic map(
            re_multiplicator=>-16364, --- -0.998779296875 + j0.0490112304688
            im_multiplicator=>803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1684),
            data_im_in=>first_stage_im_out(1684),
            product_re_out=>mul_re_out(1684),
            product_im_out=>mul_im_out(1684)
        );

    UMUL_1685 : complex_multiplier
    generic map(
            re_multiplicator=>-16028, --- -0.978271484375 + j0.207092285156
            im_multiplicator=>3393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1685),
            data_im_in=>first_stage_im_out(1685),
            product_re_out=>mul_re_out(1685),
            product_im_out=>mul_im_out(1685)
        );

    UMUL_1686 : complex_multiplier
    generic map(
            re_multiplicator=>-15286, --- -0.932983398438 + j0.35986328125
            im_multiplicator=>5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1686),
            data_im_in=>first_stage_im_out(1686),
            product_re_out=>mul_re_out(1686),
            product_im_out=>mul_im_out(1686)
        );

    UMUL_1687 : complex_multiplier
    generic map(
            re_multiplicator=>-14155, --- -0.863952636719 + j0.503479003906
            im_multiplicator=>8249
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1687),
            data_im_in=>first_stage_im_out(1687),
            product_re_out=>mul_re_out(1687),
            product_im_out=>mul_im_out(1687)
        );

    UMUL_1688 : complex_multiplier
    generic map(
            re_multiplicator=>-12665, --- -0.773010253906 + j0.634338378906
            im_multiplicator=>10393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1688),
            data_im_in=>first_stage_im_out(1688),
            product_re_out=>mul_re_out(1688),
            product_im_out=>mul_im_out(1688)
        );

    UMUL_1689 : complex_multiplier
    generic map(
            re_multiplicator=>-10853, --- -0.662414550781 + j0.749084472656
            im_multiplicator=>12273
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1689),
            data_im_in=>first_stage_im_out(1689),
            product_re_out=>mul_re_out(1689),
            product_im_out=>mul_im_out(1689)
        );

    UMUL_1690 : complex_multiplier
    generic map(
            re_multiplicator=>-8765, --- -0.534973144531 + j0.844848632812
            im_multiplicator=>13842
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1690),
            data_im_in=>first_stage_im_out(1690),
            product_re_out=>mul_re_out(1690),
            product_im_out=>mul_im_out(1690)
        );

    UMUL_1691 : complex_multiplier
    generic map(
            re_multiplicator=>-6455, --- -0.393981933594 + j0.919067382812
            im_multiplicator=>15058
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1691),
            data_im_in=>first_stage_im_out(1691),
            product_re_out=>mul_re_out(1691),
            product_im_out=>mul_im_out(1691)
        );

    UMUL_1692 : complex_multiplier
    generic map(
            re_multiplicator=>-3980, --- -0.242919921875 + j0.969970703125
            im_multiplicator=>15892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1692),
            data_im_in=>first_stage_im_out(1692),
            product_re_out=>mul_re_out(1692),
            product_im_out=>mul_im_out(1692)
        );

    UMUL_1693 : complex_multiplier
    generic map(
            re_multiplicator=>-1405, --- -0.0857543945312 + j0.996276855469
            im_multiplicator=>16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1693),
            data_im_in=>first_stage_im_out(1693),
            product_re_out=>mul_re_out(1693),
            product_im_out=>mul_im_out(1693)
        );

    UMUL_1694 : complex_multiplier
    generic map(
            re_multiplicator=>1205, --- 0.0735473632812 + j0.997253417969
            im_multiplicator=>16339
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1694),
            data_im_in=>first_stage_im_out(1694),
            product_re_out=>mul_re_out(1694),
            product_im_out=>mul_im_out(1694)
        );

    UMUL_1695 : complex_multiplier
    generic map(
            re_multiplicator=>3785, --- 0.231018066406 + j0.972900390625
            im_multiplicator=>15940
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1695),
            data_im_in=>first_stage_im_out(1695),
            product_re_out=>mul_re_out(1695),
            product_im_out=>mul_im_out(1695)
        );

    UDELAY_1696_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1696),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1696)
        );
    UDELAY_1696_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1696),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1696)
        );
    USHIFTER_1696_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1696),
            data_out=>mul_re_out(1696)
        );
    USHIFTER_1696_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1696),
            data_out=>mul_im_out(1696)
        );

    UMUL_1697 : complex_multiplier
    generic map(
            re_multiplicator=>16167, --- 0.986755371094 + j-0.161865234375
            im_multiplicator=>-2652
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1697),
            data_im_in=>first_stage_im_out(1697),
            product_re_out=>mul_re_out(1697),
            product_im_out=>mul_im_out(1697)
        );

    UMUL_1698 : complex_multiplier
    generic map(
            re_multiplicator=>15525, --- 0.947570800781 + j-0.319458007812
            im_multiplicator=>-5234
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1698),
            data_im_in=>first_stage_im_out(1698),
            product_re_out=>mul_re_out(1698),
            product_im_out=>mul_im_out(1698)
        );

    UMUL_1699 : complex_multiplier
    generic map(
            re_multiplicator=>14473, --- 0.883361816406 + j-0.468627929688
            im_multiplicator=>-7678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1699),
            data_im_in=>first_stage_im_out(1699),
            product_re_out=>mul_re_out(1699),
            product_im_out=>mul_im_out(1699)
        );

    UMUL_1700 : complex_multiplier
    generic map(
            re_multiplicator=>13038, --- 0.795776367188 + j-0.60546875
            im_multiplicator=>-9920
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1700),
            data_im_in=>first_stage_im_out(1700),
            product_re_out=>mul_re_out(1700),
            product_im_out=>mul_im_out(1700)
        );

    UMUL_1701 : complex_multiplier
    generic map(
            re_multiplicator=>11260, --- 0.687255859375 + j-0.726318359375
            im_multiplicator=>-11900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1701),
            data_im_in=>first_stage_im_out(1701),
            product_re_out=>mul_re_out(1701),
            product_im_out=>mul_im_out(1701)
        );

    UMUL_1702 : complex_multiplier
    generic map(
            re_multiplicator=>9185, --- 0.560607910156 + j-0.828002929688
            im_multiplicator=>-13566
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1702),
            data_im_in=>first_stage_im_out(1702),
            product_re_out=>mul_re_out(1702),
            product_im_out=>mul_im_out(1702)
        );

    UMUL_1703 : complex_multiplier
    generic map(
            re_multiplicator=>6868, --- 0.419189453125 + j-0.907836914062
            im_multiplicator=>-14874
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1703),
            data_im_in=>first_stage_im_out(1703),
            product_re_out=>mul_re_out(1703),
            product_im_out=>mul_im_out(1703)
        );

    UMUL_1704 : complex_multiplier
    generic map(
            re_multiplicator=>4369, --- 0.266662597656 + j-0.963745117188
            im_multiplicator=>-15790
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1704),
            data_im_in=>first_stage_im_out(1704),
            product_re_out=>mul_re_out(1704),
            product_im_out=>mul_im_out(1704)
        );

    UMUL_1705 : complex_multiplier
    generic map(
            re_multiplicator=>1755, --- 0.107116699219 + j-0.994201660156
            im_multiplicator=>-16289
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1705),
            data_im_in=>first_stage_im_out(1705),
            product_re_out=>mul_re_out(1705),
            product_im_out=>mul_im_out(1705)
        );

    UMUL_1706 : complex_multiplier
    generic map(
            re_multiplicator=>-904, --- -0.05517578125 + j-0.998474121094
            im_multiplicator=>-16359
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1706),
            data_im_in=>first_stage_im_out(1706),
            product_re_out=>mul_re_out(1706),
            product_im_out=>mul_im_out(1706)
        );

    UMUL_1707 : complex_multiplier
    generic map(
            re_multiplicator=>-3540, --- -0.216064453125 + j-0.976318359375
            im_multiplicator=>-15996
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1707),
            data_im_in=>first_stage_im_out(1707),
            product_re_out=>mul_re_out(1707),
            product_im_out=>mul_im_out(1707)
        );

    UMUL_1708 : complex_multiplier
    generic map(
            re_multiplicator=>-6083, --- -0.371276855469 + j-0.928466796875
            im_multiplicator=>-15212
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1708),
            data_im_in=>first_stage_im_out(1708),
            product_re_out=>mul_re_out(1708),
            product_im_out=>mul_im_out(1708)
        );

    UMUL_1709 : complex_multiplier
    generic map(
            re_multiplicator=>-8466, --- -0.516723632812 + j-0.856140136719
            im_multiplicator=>-14027
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1709),
            data_im_in=>first_stage_im_out(1709),
            product_re_out=>mul_re_out(1709),
            product_im_out=>mul_im_out(1709)
        );

    UMUL_1710 : complex_multiplier
    generic map(
            re_multiplicator=>-10625, --- -0.648498535156 + j-0.761169433594
            im_multiplicator=>-12471
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1710),
            data_im_in=>first_stage_im_out(1710),
            product_re_out=>mul_re_out(1710),
            product_im_out=>mul_im_out(1710)
        );

    UMUL_1711 : complex_multiplier
    generic map(
            re_multiplicator=>-12504, --- -0.76318359375 + j-0.646118164062
            im_multiplicator=>-10586
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1711),
            data_im_in=>first_stage_im_out(1711),
            product_re_out=>mul_re_out(1711),
            product_im_out=>mul_im_out(1711)
        );

    UMUL_1712 : complex_multiplier
    generic map(
            re_multiplicator=>-14053, --- -0.857727050781 + j-0.514099121094
            im_multiplicator=>-8423
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1712),
            data_im_in=>first_stage_im_out(1712),
            product_re_out=>mul_re_out(1712),
            product_im_out=>mul_im_out(1712)
        );

    UMUL_1713 : complex_multiplier
    generic map(
            re_multiplicator=>-15231, --- -0.929626464844 + j-0.368408203125
            im_multiplicator=>-6036
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1713),
            data_im_in=>first_stage_im_out(1713),
            product_re_out=>mul_re_out(1713),
            product_im_out=>mul_im_out(1713)
        );

    UMUL_1714 : complex_multiplier
    generic map(
            re_multiplicator=>-16007, --- -0.976989746094 + j-0.213073730469
            im_multiplicator=>-3491
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1714),
            data_im_in=>first_stage_im_out(1714),
            product_re_out=>mul_re_out(1714),
            product_im_out=>mul_im_out(1714)
        );

    UMUL_1715 : complex_multiplier
    generic map(
            re_multiplicator=>-16361, --- -0.998596191406 + j-0.0521240234375
            im_multiplicator=>-854
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1715),
            data_im_in=>first_stage_im_out(1715),
            product_re_out=>mul_re_out(1715),
            product_im_out=>mul_im_out(1715)
        );

    UMUL_1716 : complex_multiplier
    generic map(
            re_multiplicator=>-16284, --- -0.993896484375 + j0.110168457031
            im_multiplicator=>1805
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1716),
            data_im_in=>first_stage_im_out(1716),
            product_re_out=>mul_re_out(1716),
            product_im_out=>mul_im_out(1716)
        );

    UMUL_1717 : complex_multiplier
    generic map(
            re_multiplicator=>-15777, --- -0.962951660156 + j0.269653320312
            im_multiplicator=>4418
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1717),
            data_im_in=>first_stage_im_out(1717),
            product_re_out=>mul_re_out(1717),
            product_im_out=>mul_im_out(1717)
        );

    UMUL_1718 : complex_multiplier
    generic map(
            re_multiplicator=>-14853, --- -0.906555175781 + j0.421997070312
            im_multiplicator=>6914
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1718),
            data_im_in=>first_stage_im_out(1718),
            product_re_out=>mul_re_out(1718),
            product_im_out=>mul_im_out(1718)
        );

    UMUL_1719 : complex_multiplier
    generic map(
            re_multiplicator=>-13538, --- -0.826293945312 + j0.563171386719
            im_multiplicator=>9227
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1719),
            data_im_in=>first_stage_im_out(1719),
            product_re_out=>mul_re_out(1719),
            product_im_out=>mul_im_out(1719)
        );

    UMUL_1720 : complex_multiplier
    generic map(
            re_multiplicator=>-11866, --- -0.724243164062 + j0.689514160156
            im_multiplicator=>11297
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1720),
            data_im_in=>first_stage_im_out(1720),
            product_re_out=>mul_re_out(1720),
            product_im_out=>mul_im_out(1720)
        );

    UMUL_1721 : complex_multiplier
    generic map(
            re_multiplicator=>-9880, --- -0.60302734375 + j0.797668457031
            im_multiplicator=>13069
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1721),
            data_im_in=>first_stage_im_out(1721),
            product_re_out=>mul_re_out(1721),
            product_im_out=>mul_im_out(1721)
        );

    UMUL_1722 : complex_multiplier
    generic map(
            re_multiplicator=>-7634, --- -0.465942382812 + j0.884765625
            im_multiplicator=>14496
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1722),
            data_im_in=>first_stage_im_out(1722),
            product_re_out=>mul_re_out(1722),
            product_im_out=>mul_im_out(1722)
        );

    UMUL_1723 : complex_multiplier
    generic map(
            re_multiplicator=>-5187, --- -0.316589355469 + j0.948547363281
            im_multiplicator=>15541
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1723),
            data_im_in=>first_stage_im_out(1723),
            product_re_out=>mul_re_out(1723),
            product_im_out=>mul_im_out(1723)
        );

    UMUL_1724 : complex_multiplier
    generic map(
            re_multiplicator=>-2602, --- -0.158813476562 + j0.987243652344
            im_multiplicator=>16175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1724),
            data_im_in=>first_stage_im_out(1724),
            product_re_out=>mul_re_out(1724),
            product_im_out=>mul_im_out(1724)
        );

    UMUL_1725 : complex_multiplier
    generic map(
            re_multiplicator=>50, --- 0.0030517578125 + j0.999938964844
            im_multiplicator=>16383
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1725),
            data_im_in=>first_stage_im_out(1725),
            product_re_out=>mul_re_out(1725),
            product_im_out=>mul_im_out(1725)
        );

    UMUL_1726 : complex_multiplier
    generic map(
            re_multiplicator=>2701, --- 0.164855957031 + j0.986267089844
            im_multiplicator=>16159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1726),
            data_im_in=>first_stage_im_out(1726),
            product_re_out=>mul_re_out(1726),
            product_im_out=>mul_im_out(1726)
        );

    UMUL_1727 : complex_multiplier
    generic map(
            re_multiplicator=>5282, --- 0.322387695312 + j0.946594238281
            im_multiplicator=>15509
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1727),
            data_im_in=>first_stage_im_out(1727),
            product_re_out=>mul_re_out(1727),
            product_im_out=>mul_im_out(1727)
        );

    UDELAY_1728_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1728),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1728)
        );
    UDELAY_1728_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1728),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1728)
        );
    USHIFTER_1728_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1728),
            data_out=>mul_re_out(1728)
        );
    USHIFTER_1728_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1728),
            data_out=>mul_im_out(1728)
        );

    UMUL_1729 : complex_multiplier
    generic map(
            re_multiplicator=>16159, --- 0.986267089844 + j-0.164855957031
            im_multiplicator=>-2701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1729),
            data_im_in=>first_stage_im_out(1729),
            product_re_out=>mul_re_out(1729),
            product_im_out=>mul_im_out(1729)
        );

    UMUL_1730 : complex_multiplier
    generic map(
            re_multiplicator=>15492, --- 0.945556640625 + j-0.325256347656
            im_multiplicator=>-5329
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1730),
            data_im_in=>first_stage_im_out(1730),
            product_re_out=>mul_re_out(1730),
            product_im_out=>mul_im_out(1730)
        );

    UMUL_1731 : complex_multiplier
    generic map(
            re_multiplicator=>14401, --- 0.878967285156 + j-0.476745605469
            im_multiplicator=>-7811
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1731),
            data_im_in=>first_stage_im_out(1731),
            product_re_out=>mul_re_out(1731),
            product_im_out=>mul_im_out(1731)
        );

    UMUL_1732 : complex_multiplier
    generic map(
            re_multiplicator=>12916, --- 0.788330078125 + j-0.615173339844
            im_multiplicator=>-10079
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1732),
            data_im_in=>first_stage_im_out(1732),
            product_re_out=>mul_re_out(1732),
            product_im_out=>mul_im_out(1732)
        );

    UMUL_1733 : complex_multiplier
    generic map(
            re_multiplicator=>11077, --- 0.676086425781 + j-0.73681640625
            im_multiplicator=>-12072
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1733),
            data_im_in=>first_stage_im_out(1733),
            product_re_out=>mul_re_out(1733),
            product_im_out=>mul_im_out(1733)
        );

    UMUL_1734 : complex_multiplier
    generic map(
            re_multiplicator=>8934, --- 0.545288085938 + j-0.838195800781
            im_multiplicator=>-13733
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1734),
            data_im_in=>first_stage_im_out(1734),
            product_re_out=>mul_re_out(1734),
            product_im_out=>mul_im_out(1734)
        );

    UMUL_1735 : complex_multiplier
    generic map(
            re_multiplicator=>6547, --- 0.399597167969 + j-0.916625976562
            im_multiplicator=>-15018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1735),
            data_im_in=>first_stage_im_out(1735),
            product_re_out=>mul_re_out(1735),
            product_im_out=>mul_im_out(1735)
        );

    UMUL_1736 : complex_multiplier
    generic map(
            re_multiplicator=>3980, --- 0.242919921875 + j-0.969970703125
            im_multiplicator=>-15892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1736),
            data_im_in=>first_stage_im_out(1736),
            product_re_out=>mul_re_out(1736),
            product_im_out=>mul_im_out(1736)
        );

    UMUL_1737 : complex_multiplier
    generic map(
            re_multiplicator=>1305, --- 0.0796508789062 + j-0.996765136719
            im_multiplicator=>-16331
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1737),
            data_im_in=>first_stage_im_out(1737),
            product_re_out=>mul_re_out(1737),
            product_im_out=>mul_im_out(1737)
        );

    UMUL_1738 : complex_multiplier
    generic map(
            re_multiplicator=>-1405, --- -0.0857543945312 + j-0.996276855469
            im_multiplicator=>-16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1738),
            data_im_in=>first_stage_im_out(1738),
            product_re_out=>mul_re_out(1738),
            product_im_out=>mul_im_out(1738)
        );

    UMUL_1739 : complex_multiplier
    generic map(
            re_multiplicator=>-4078, --- -0.248901367188 + j-0.968505859375
            im_multiplicator=>-15868
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1739),
            data_im_in=>first_stage_im_out(1739),
            product_re_out=>mul_re_out(1739),
            product_im_out=>mul_im_out(1739)
        );

    UMUL_1740 : complex_multiplier
    generic map(
            re_multiplicator=>-6639, --- -0.405212402344 + j-0.914184570312
            im_multiplicator=>-14978
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1740),
            data_im_in=>first_stage_im_out(1740),
            product_re_out=>mul_re_out(1740),
            product_im_out=>mul_im_out(1740)
        );

    UMUL_1741 : complex_multiplier
    generic map(
            re_multiplicator=>-9018, --- -0.550415039062 + j-0.834838867188
            im_multiplicator=>-13678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1741),
            data_im_in=>first_stage_im_out(1741),
            product_re_out=>mul_re_out(1741),
            product_im_out=>mul_im_out(1741)
        );

    UMUL_1742 : complex_multiplier
    generic map(
            re_multiplicator=>-11150, --- -0.680541992188 + j-0.732604980469
            im_multiplicator=>-12003
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1742),
            data_im_in=>first_stage_im_out(1742),
            product_re_out=>mul_re_out(1742),
            product_im_out=>mul_im_out(1742)
        );

    UMUL_1743 : complex_multiplier
    generic map(
            re_multiplicator=>-12977, --- -0.792053222656 + j-0.6103515625
            im_multiplicator=>-10000
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1743),
            data_im_in=>first_stage_im_out(1743),
            product_re_out=>mul_re_out(1743),
            product_im_out=>mul_im_out(1743)
        );

    UMUL_1744 : complex_multiplier
    generic map(
            re_multiplicator=>-14449, --- -0.881896972656 + j-0.471374511719
            im_multiplicator=>-7723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1744),
            data_im_in=>first_stage_im_out(1744),
            product_re_out=>mul_re_out(1744),
            product_im_out=>mul_im_out(1744)
        );

    UMUL_1745 : complex_multiplier
    generic map(
            re_multiplicator=>-15525, --- -0.947570800781 + j-0.319458007812
            im_multiplicator=>-5234
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1745),
            data_im_in=>first_stage_im_out(1745),
            product_re_out=>mul_re_out(1745),
            product_im_out=>mul_im_out(1745)
        );

    UMUL_1746 : complex_multiplier
    generic map(
            re_multiplicator=>-16175, --- -0.987243652344 + j-0.158813476562
            im_multiplicator=>-2602
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1746),
            data_im_in=>first_stage_im_out(1746),
            product_re_out=>mul_re_out(1746),
            product_im_out=>mul_im_out(1746)
        );

    UMUL_1747 : complex_multiplier
    generic map(
            re_multiplicator=>-16383, --- -0.999938964844 + j0.006103515625
            im_multiplicator=>100
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1747),
            data_im_in=>first_stage_im_out(1747),
            product_re_out=>mul_re_out(1747),
            product_im_out=>mul_im_out(1747)
        );

    UMUL_1748 : complex_multiplier
    generic map(
            re_multiplicator=>-16142, --- -0.985229492188 + j0.170959472656
            im_multiplicator=>2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1748),
            data_im_in=>first_stage_im_out(1748),
            product_re_out=>mul_re_out(1748),
            product_im_out=>mul_im_out(1748)
        );

    UMUL_1749 : complex_multiplier
    generic map(
            re_multiplicator=>-15459, --- -0.943542480469 + j0.3310546875
            im_multiplicator=>5424
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1749),
            data_im_in=>first_stage_im_out(1749),
            product_re_out=>mul_re_out(1749),
            product_im_out=>mul_im_out(1749)
        );

    UMUL_1750 : complex_multiplier
    generic map(
            re_multiplicator=>-14353, --- -0.876037597656 + j0.482177734375
            im_multiplicator=>7900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1750),
            data_im_in=>first_stage_im_out(1750),
            product_re_out=>mul_re_out(1750),
            product_im_out=>mul_im_out(1750)
        );

    UMUL_1751 : complex_multiplier
    generic map(
            re_multiplicator=>-12854, --- -0.784545898438 + j0.620056152344
            im_multiplicator=>10159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1751),
            data_im_in=>first_stage_im_out(1751),
            product_re_out=>mul_re_out(1751),
            product_im_out=>mul_im_out(1751)
        );

    UMUL_1752 : complex_multiplier
    generic map(
            re_multiplicator=>-11002, --- -0.671508789062 + j0.740905761719
            im_multiplicator=>12139
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1752),
            data_im_in=>first_stage_im_out(1752),
            product_re_out=>mul_re_out(1752),
            product_im_out=>mul_im_out(1752)
        );

    UMUL_1753 : complex_multiplier
    generic map(
            re_multiplicator=>-8850, --- -0.540161132812 + j0.841552734375
            im_multiplicator=>13788
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1753),
            data_im_in=>first_stage_im_out(1753),
            product_re_out=>mul_re_out(1753),
            product_im_out=>mul_im_out(1753)
        );

    UMUL_1754 : complex_multiplier
    generic map(
            re_multiplicator=>-6455, --- -0.393981933594 + j0.919067382812
            im_multiplicator=>15058
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1754),
            data_im_in=>first_stage_im_out(1754),
            product_re_out=>mul_re_out(1754),
            product_im_out=>mul_im_out(1754)
        );

    UMUL_1755 : complex_multiplier
    generic map(
            re_multiplicator=>-3883, --- -0.236999511719 + j0.971496582031
            im_multiplicator=>15917
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1755),
            data_im_in=>first_stage_im_out(1755),
            product_re_out=>mul_re_out(1755),
            product_im_out=>mul_im_out(1755)
        );

    UMUL_1756 : complex_multiplier
    generic map(
            re_multiplicator=>-1205, --- -0.0735473632812 + j0.997253417969
            im_multiplicator=>16339
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1756),
            data_im_in=>first_stage_im_out(1756),
            product_re_out=>mul_re_out(1756),
            product_im_out=>mul_im_out(1756)
        );

    UMUL_1757 : complex_multiplier
    generic map(
            re_multiplicator=>1505, --- 0.0918579101562 + j0.995727539062
            im_multiplicator=>16314
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1757),
            data_im_in=>first_stage_im_out(1757),
            product_re_out=>mul_re_out(1757),
            product_im_out=>mul_im_out(1757)
        );

    UMUL_1758 : complex_multiplier
    generic map(
            re_multiplicator=>4175, --- 0.254821777344 + j0.966918945312
            im_multiplicator=>15842
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1758),
            data_im_in=>first_stage_im_out(1758),
            product_re_out=>mul_re_out(1758),
            product_im_out=>mul_im_out(1758)
        );

    UMUL_1759 : complex_multiplier
    generic map(
            re_multiplicator=>6731, --- 0.410827636719 + j0.911682128906
            im_multiplicator=>14937
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1759),
            data_im_in=>first_stage_im_out(1759),
            product_re_out=>mul_re_out(1759),
            product_im_out=>mul_im_out(1759)
        );

    UDELAY_1760_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1760),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1760)
        );
    UDELAY_1760_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1760),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1760)
        );
    USHIFTER_1760_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1760),
            data_out=>mul_re_out(1760)
        );
    USHIFTER_1760_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1760),
            data_out=>mul_im_out(1760)
        );

    UMUL_1761 : complex_multiplier
    generic map(
            re_multiplicator=>16151, --- 0.985778808594 + j-0.167907714844
            im_multiplicator=>-2751
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1761),
            data_im_in=>first_stage_im_out(1761),
            product_re_out=>mul_re_out(1761),
            product_im_out=>mul_im_out(1761)
        );

    UMUL_1762 : complex_multiplier
    generic map(
            re_multiplicator=>15459, --- 0.943542480469 + j-0.3310546875
            im_multiplicator=>-5424
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1762),
            data_im_in=>first_stage_im_out(1762),
            product_re_out=>mul_re_out(1762),
            product_im_out=>mul_im_out(1762)
        );

    UMUL_1763 : complex_multiplier
    generic map(
            re_multiplicator=>14329, --- 0.874572753906 + j-0.48486328125
            im_multiplicator=>-7944
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1763),
            data_im_in=>first_stage_im_out(1763),
            product_re_out=>mul_re_out(1763),
            product_im_out=>mul_im_out(1763)
        );

    UMUL_1764 : complex_multiplier
    generic map(
            re_multiplicator=>12791, --- 0.780700683594 + j-0.624816894531
            im_multiplicator=>-10237
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1764),
            data_im_in=>first_stage_im_out(1764),
            product_re_out=>mul_re_out(1764),
            product_im_out=>mul_im_out(1764)
        );

    UMUL_1765 : complex_multiplier
    generic map(
            re_multiplicator=>10890, --- 0.664672851562 + j-0.7470703125
            im_multiplicator=>-12240
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1765),
            data_im_in=>first_stage_im_out(1765),
            product_re_out=>mul_re_out(1765),
            product_im_out=>mul_im_out(1765)
        );

    UMUL_1766 : complex_multiplier
    generic map(
            re_multiplicator=>8680, --- 0.52978515625 + j-0.848083496094
            im_multiplicator=>-13895
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1766),
            data_im_in=>first_stage_im_out(1766),
            product_re_out=>mul_re_out(1766),
            product_im_out=>mul_im_out(1766)
        );

    UMUL_1767 : complex_multiplier
    generic map(
            re_multiplicator=>6223, --- 0.379821777344 + j-0.925048828125
            im_multiplicator=>-15156
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1767),
            data_im_in=>first_stage_im_out(1767),
            product_re_out=>mul_re_out(1767),
            product_im_out=>mul_im_out(1767)
        );

    UMUL_1768 : complex_multiplier
    generic map(
            re_multiplicator=>3589, --- 0.219055175781 + j-0.975646972656
            im_multiplicator=>-15985
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1768),
            data_im_in=>first_stage_im_out(1768),
            product_re_out=>mul_re_out(1768),
            product_im_out=>mul_im_out(1768)
        );

    UMUL_1769 : complex_multiplier
    generic map(
            re_multiplicator=>854, --- 0.0521240234375 + j-0.998596191406
            im_multiplicator=>-16361
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1769),
            data_im_in=>first_stage_im_out(1769),
            product_re_out=>mul_re_out(1769),
            product_im_out=>mul_im_out(1769)
        );

    UMUL_1770 : complex_multiplier
    generic map(
            re_multiplicator=>-1905, --- -0.116271972656 + j-0.9931640625
            im_multiplicator=>-16272
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1770),
            data_im_in=>first_stage_im_out(1770),
            product_re_out=>mul_re_out(1770),
            product_im_out=>mul_im_out(1770)
        );

    UMUL_1771 : complex_multiplier
    generic map(
            re_multiplicator=>-4611, --- -0.281433105469 + j-0.959533691406
            im_multiplicator=>-15721
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1771),
            data_im_in=>first_stage_im_out(1771),
            product_re_out=>mul_re_out(1771),
            product_im_out=>mul_im_out(1771)
        );

    UMUL_1772 : complex_multiplier
    generic map(
            re_multiplicator=>-7186, --- -0.438598632812 + j-0.898620605469
            im_multiplicator=>-14723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1772),
            data_im_in=>first_stage_im_out(1772),
            product_re_out=>mul_re_out(1772),
            product_im_out=>mul_im_out(1772)
        );

    UMUL_1773 : complex_multiplier
    generic map(
            re_multiplicator=>-9556, --- -0.583251953125 + j-0.812194824219
            im_multiplicator=>-13307
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1773),
            data_im_in=>first_stage_im_out(1773),
            product_re_out=>mul_re_out(1773),
            product_im_out=>mul_im_out(1773)
        );

    UMUL_1774 : complex_multiplier
    generic map(
            re_multiplicator=>-11656, --- -0.71142578125 + j-0.702697753906
            im_multiplicator=>-11513
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1774),
            data_im_in=>first_stage_im_out(1774),
            product_re_out=>mul_re_out(1774),
            product_im_out=>mul_im_out(1774)
        );

    UMUL_1775 : complex_multiplier
    generic map(
            re_multiplicator=>-13424, --- -0.8193359375 + j-0.5732421875
            im_multiplicator=>-9392
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1775),
            data_im_in=>first_stage_im_out(1775),
            product_re_out=>mul_re_out(1775),
            product_im_out=>mul_im_out(1775)
        );

    UMUL_1776 : complex_multiplier
    generic map(
            re_multiplicator=>-14810, --- -0.903930664062 + j-0.427551269531
            im_multiplicator=>-7005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1776),
            data_im_in=>first_stage_im_out(1776),
            product_re_out=>mul_re_out(1776),
            product_im_out=>mul_im_out(1776)
        );

    UMUL_1777 : complex_multiplier
    generic map(
            re_multiplicator=>-15777, --- -0.962951660156 + j-0.269653320312
            im_multiplicator=>-4418
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1777),
            data_im_in=>first_stage_im_out(1777),
            product_re_out=>mul_re_out(1777),
            product_im_out=>mul_im_out(1777)
        );

    UMUL_1778 : complex_multiplier
    generic map(
            re_multiplicator=>-16294, --- -0.994506835938 + j-0.104064941406
            im_multiplicator=>-1705
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1778),
            data_im_in=>first_stage_im_out(1778),
            product_re_out=>mul_re_out(1778),
            product_im_out=>mul_im_out(1778)
        );

    UMUL_1779 : complex_multiplier
    generic map(
            re_multiplicator=>-16350, --- -0.997924804688 + j0.0643310546875
            im_multiplicator=>1054
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1779),
            data_im_in=>first_stage_im_out(1779),
            product_re_out=>mul_re_out(1779),
            product_im_out=>mul_im_out(1779)
        );

    UMUL_1780 : complex_multiplier
    generic map(
            re_multiplicator=>-15940, --- -0.972900390625 + j0.231018066406
            im_multiplicator=>3785
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1780),
            data_im_in=>first_stage_im_out(1780),
            product_re_out=>mul_re_out(1780),
            product_im_out=>mul_im_out(1780)
        );

    UMUL_1781 : complex_multiplier
    generic map(
            re_multiplicator=>-15078, --- -0.920288085938 + j0.39111328125
            im_multiplicator=>6408
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1781),
            data_im_in=>first_stage_im_out(1781),
            product_re_out=>mul_re_out(1781),
            product_im_out=>mul_im_out(1781)
        );

    UMUL_1782 : complex_multiplier
    generic map(
            re_multiplicator=>-13788, --- -0.841552734375 + j0.540161132812
            im_multiplicator=>8850
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1782),
            data_im_in=>first_stage_im_out(1782),
            product_re_out=>mul_re_out(1782),
            product_im_out=>mul_im_out(1782)
        );

    UMUL_1783 : complex_multiplier
    generic map(
            re_multiplicator=>-12105, --- -0.738830566406 + j0.673828125
            im_multiplicator=>11040
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1783),
            data_im_in=>first_stage_im_out(1783),
            product_re_out=>mul_re_out(1783),
            product_im_out=>mul_im_out(1783)
        );

    UMUL_1784 : complex_multiplier
    generic map(
            re_multiplicator=>-10079, --- -0.615173339844 + j0.788330078125
            im_multiplicator=>12916
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1784),
            data_im_in=>first_stage_im_out(1784),
            product_re_out=>mul_re_out(1784),
            product_im_out=>mul_im_out(1784)
        );

    UMUL_1785 : complex_multiplier
    generic map(
            re_multiplicator=>-7767, --- -0.474060058594 + j0.880432128906
            im_multiplicator=>14425
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1785),
            data_im_in=>first_stage_im_out(1785),
            product_re_out=>mul_re_out(1785),
            product_im_out=>mul_im_out(1785)
        );

    UMUL_1786 : complex_multiplier
    generic map(
            re_multiplicator=>-5234, --- -0.319458007812 + j0.947570800781
            im_multiplicator=>15525
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1786),
            data_im_in=>first_stage_im_out(1786),
            product_re_out=>mul_re_out(1786),
            product_im_out=>mul_im_out(1786)
        );

    UMUL_1787 : complex_multiplier
    generic map(
            re_multiplicator=>-2553, --- -0.155822753906 + j0.987731933594
            im_multiplicator=>16183
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1787),
            data_im_in=>first_stage_im_out(1787),
            product_re_out=>mul_re_out(1787),
            product_im_out=>mul_im_out(1787)
        );

    UMUL_1788 : complex_multiplier
    generic map(
            re_multiplicator=>201, --- 0.0122680664062 + j0.999877929688
            im_multiplicator=>16382
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1788),
            data_im_in=>first_stage_im_out(1788),
            product_re_out=>mul_re_out(1788),
            product_im_out=>mul_im_out(1788)
        );

    UMUL_1789 : complex_multiplier
    generic map(
            re_multiplicator=>2949, --- 0.179992675781 + j0.983642578125
            im_multiplicator=>16116
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1789),
            data_im_in=>first_stage_im_out(1789),
            product_re_out=>mul_re_out(1789),
            product_im_out=>mul_im_out(1789)
        );

    UMUL_1790 : complex_multiplier
    generic map(
            re_multiplicator=>5614, --- 0.342651367188 + j0.939453125
            im_multiplicator=>15392
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1790),
            data_im_in=>first_stage_im_out(1790),
            product_re_out=>mul_re_out(1790),
            product_im_out=>mul_im_out(1790)
        );

    UMUL_1791 : complex_multiplier
    generic map(
            re_multiplicator=>8119, --- 0.495544433594 + j0.868530273438
            im_multiplicator=>14230
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1791),
            data_im_in=>first_stage_im_out(1791),
            product_re_out=>mul_re_out(1791),
            product_im_out=>mul_im_out(1791)
        );

    UDELAY_1792_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1792),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1792)
        );
    UDELAY_1792_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1792),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1792)
        );
    USHIFTER_1792_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1792),
            data_out=>mul_re_out(1792)
        );
    USHIFTER_1792_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1792),
            data_out=>mul_im_out(1792)
        );

    UMUL_1793 : complex_multiplier
    generic map(
            re_multiplicator=>16142, --- 0.985229492188 + j-0.170959472656
            im_multiplicator=>-2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1793),
            data_im_in=>first_stage_im_out(1793),
            product_re_out=>mul_re_out(1793),
            product_im_out=>mul_im_out(1793)
        );

    UMUL_1794 : complex_multiplier
    generic map(
            re_multiplicator=>15426, --- 0.941528320312 + j-0.336853027344
            im_multiplicator=>-5519
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1794),
            data_im_in=>first_stage_im_out(1794),
            product_re_out=>mul_re_out(1794),
            product_im_out=>mul_im_out(1794)
        );

    UMUL_1795 : complex_multiplier
    generic map(
            re_multiplicator=>14255, --- 0.870056152344 + j-0.492858886719
            im_multiplicator=>-8075
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1795),
            data_im_in=>first_stage_im_out(1795),
            product_re_out=>mul_re_out(1795),
            product_im_out=>mul_im_out(1795)
        );

    UMUL_1796 : complex_multiplier
    generic map(
            re_multiplicator=>12665, --- 0.773010253906 + j-0.634338378906
            im_multiplicator=>-10393
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1796),
            data_im_in=>first_stage_im_out(1796),
            product_re_out=>mul_re_out(1796),
            product_im_out=>mul_im_out(1796)
        );

    UMUL_1797 : complex_multiplier
    generic map(
            re_multiplicator=>10701, --- 0.653137207031 + j-0.757202148438
            im_multiplicator=>-12406
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1797),
            data_im_in=>first_stage_im_out(1797),
            product_re_out=>mul_re_out(1797),
            product_im_out=>mul_im_out(1797)
        );

    UMUL_1798 : complex_multiplier
    generic map(
            re_multiplicator=>8423, --- 0.514099121094 + j-0.857727050781
            im_multiplicator=>-14053
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1798),
            data_im_in=>first_stage_im_out(1798),
            product_re_out=>mul_re_out(1798),
            product_im_out=>mul_im_out(1798)
        );

    UMUL_1799 : complex_multiplier
    generic map(
            re_multiplicator=>5896, --- 0.35986328125 + j-0.932983398438
            im_multiplicator=>-15286
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1799),
            data_im_in=>first_stage_im_out(1799),
            product_re_out=>mul_re_out(1799),
            product_im_out=>mul_im_out(1799)
        );

    UMUL_1800 : complex_multiplier
    generic map(
            re_multiplicator=>3196, --- 0.195068359375 + j-0.980773925781
            im_multiplicator=>-16069
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1800),
            data_im_in=>first_stage_im_out(1800),
            product_re_out=>mul_re_out(1800),
            product_im_out=>mul_im_out(1800)
        );

    UMUL_1801 : complex_multiplier
    generic map(
            re_multiplicator=>402, --- 0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1801),
            data_im_in=>first_stage_im_out(1801),
            product_re_out=>mul_re_out(1801),
            product_im_out=>mul_im_out(1801)
        );

    UMUL_1802 : complex_multiplier
    generic map(
            re_multiplicator=>-2404, --- -0.146728515625 + j-0.989135742188
            im_multiplicator=>-16206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1802),
            data_im_in=>first_stage_im_out(1802),
            product_re_out=>mul_re_out(1802),
            product_im_out=>mul_im_out(1802)
        );

    UMUL_1803 : complex_multiplier
    generic map(
            re_multiplicator=>-5139, --- -0.313659667969 + j-0.949523925781
            im_multiplicator=>-15557
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1803),
            data_im_in=>first_stage_im_out(1803),
            product_re_out=>mul_re_out(1803),
            product_im_out=>mul_im_out(1803)
        );

    UMUL_1804 : complex_multiplier
    generic map(
            re_multiplicator=>-7723, --- -0.471374511719 + j-0.881896972656
            im_multiplicator=>-14449
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1804),
            data_im_in=>first_stage_im_out(1804),
            product_re_out=>mul_re_out(1804),
            product_im_out=>mul_im_out(1804)
        );

    UMUL_1805 : complex_multiplier
    generic map(
            re_multiplicator=>-10079, --- -0.615173339844 + j-0.788330078125
            im_multiplicator=>-12916
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1805),
            data_im_in=>first_stage_im_out(1805),
            product_re_out=>mul_re_out(1805),
            product_im_out=>mul_im_out(1805)
        );

    UMUL_1806 : complex_multiplier
    generic map(
            re_multiplicator=>-12139, --- -0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1806),
            data_im_in=>first_stage_im_out(1806),
            product_re_out=>mul_re_out(1806),
            product_im_out=>mul_im_out(1806)
        );

    UMUL_1807 : complex_multiplier
    generic map(
            re_multiplicator=>-13842, --- -0.844848632812 + j-0.534973144531
            im_multiplicator=>-8765
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1807),
            data_im_in=>first_stage_im_out(1807),
            product_re_out=>mul_re_out(1807),
            product_im_out=>mul_im_out(1807)
        );

    UMUL_1808 : complex_multiplier
    generic map(
            re_multiplicator=>-15136, --- -0.923828125 + j-0.382629394531
            im_multiplicator=>-6269
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1808),
            data_im_in=>first_stage_im_out(1808),
            product_re_out=>mul_re_out(1808),
            product_im_out=>mul_im_out(1808)
        );

    UMUL_1809 : complex_multiplier
    generic map(
            re_multiplicator=>-15985, --- -0.975646972656 + j-0.219055175781
            im_multiplicator=>-3589
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1809),
            data_im_in=>first_stage_im_out(1809),
            product_re_out=>mul_re_out(1809),
            product_im_out=>mul_im_out(1809)
        );

    UMUL_1810 : complex_multiplier
    generic map(
            re_multiplicator=>-16364, --- -0.998779296875 + j-0.0490112304688
            im_multiplicator=>-803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1810),
            data_im_in=>first_stage_im_out(1810),
            product_re_out=>mul_re_out(1810),
            product_im_out=>mul_im_out(1810)
        );

    UMUL_1811 : complex_multiplier
    generic map(
            re_multiplicator=>-16260, --- -0.992431640625 + j0.122375488281
            im_multiplicator=>2005
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1811),
            data_im_in=>first_stage_im_out(1811),
            product_re_out=>mul_re_out(1811),
            product_im_out=>mul_im_out(1811)
        );

    UMUL_1812 : complex_multiplier
    generic map(
            re_multiplicator=>-15678, --- -0.956909179688 + j0.290283203125
            im_multiplicator=>4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1812),
            data_im_in=>first_stage_im_out(1812),
            product_re_out=>mul_re_out(1812),
            product_im_out=>mul_im_out(1812)
        );

    UMUL_1813 : complex_multiplier
    generic map(
            re_multiplicator=>-14634, --- -0.893188476562 + j0.449584960938
            im_multiplicator=>7366
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1813),
            data_im_in=>first_stage_im_out(1813),
            product_re_out=>mul_re_out(1813),
            product_im_out=>mul_im_out(1813)
        );

    UMUL_1814 : complex_multiplier
    generic map(
            re_multiplicator=>-13159, --- -0.803161621094 + j0.595642089844
            im_multiplicator=>9759
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1814),
            data_im_in=>first_stage_im_out(1814),
            product_re_out=>mul_re_out(1814),
            product_im_out=>mul_im_out(1814)
        );

    UMUL_1815 : complex_multiplier
    generic map(
            re_multiplicator=>-11297, --- -0.689514160156 + j0.724243164062
            im_multiplicator=>11866
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1815),
            data_im_in=>first_stage_im_out(1815),
            product_re_out=>mul_re_out(1815),
            product_im_out=>mul_im_out(1815)
        );

    UMUL_1816 : complex_multiplier
    generic map(
            re_multiplicator=>-9102, --- -0.555541992188 + j0.831420898438
            im_multiplicator=>13622
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1816),
            data_im_in=>first_stage_im_out(1816),
            product_re_out=>mul_re_out(1816),
            product_im_out=>mul_im_out(1816)
        );

    UMUL_1817 : complex_multiplier
    generic map(
            re_multiplicator=>-6639, --- -0.405212402344 + j0.914184570312
            im_multiplicator=>14978
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1817),
            data_im_in=>first_stage_im_out(1817),
            product_re_out=>mul_re_out(1817),
            product_im_out=>mul_im_out(1817)
        );

    UMUL_1818 : complex_multiplier
    generic map(
            re_multiplicator=>-3980, --- -0.242919921875 + j0.969970703125
            im_multiplicator=>15892
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1818),
            data_im_in=>first_stage_im_out(1818),
            product_re_out=>mul_re_out(1818),
            product_im_out=>mul_im_out(1818)
        );

    UMUL_1819 : complex_multiplier
    generic map(
            re_multiplicator=>-1205, --- -0.0735473632812 + j0.997253417969
            im_multiplicator=>16339
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1819),
            data_im_in=>first_stage_im_out(1819),
            product_re_out=>mul_re_out(1819),
            product_im_out=>mul_im_out(1819)
        );

    UMUL_1820 : complex_multiplier
    generic map(
            re_multiplicator=>1605, --- 0.0979614257812 + j0.995178222656
            im_multiplicator=>16305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1820),
            data_im_in=>first_stage_im_out(1820),
            product_re_out=>mul_re_out(1820),
            product_im_out=>mul_im_out(1820)
        );

    UMUL_1821 : complex_multiplier
    generic map(
            re_multiplicator=>4369, --- 0.266662597656 + j0.963745117188
            im_multiplicator=>15790
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1821),
            data_im_in=>first_stage_im_out(1821),
            product_re_out=>mul_re_out(1821),
            product_im_out=>mul_im_out(1821)
        );

    UMUL_1822 : complex_multiplier
    generic map(
            re_multiplicator=>7005, --- 0.427551269531 + j0.903930664062
            im_multiplicator=>14810
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1822),
            data_im_in=>first_stage_im_out(1822),
            product_re_out=>mul_re_out(1822),
            product_im_out=>mul_im_out(1822)
        );

    UMUL_1823 : complex_multiplier
    generic map(
            re_multiplicator=>9434, --- 0.575805664062 + j0.817565917969
            im_multiplicator=>13395
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1823),
            data_im_in=>first_stage_im_out(1823),
            product_re_out=>mul_re_out(1823),
            product_im_out=>mul_im_out(1823)
        );

    UDELAY_1824_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1824),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1824)
        );
    UDELAY_1824_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1824),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1824)
        );
    USHIFTER_1824_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1824),
            data_out=>mul_re_out(1824)
        );
    USHIFTER_1824_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1824),
            data_out=>mul_im_out(1824)
        );

    UMUL_1825 : complex_multiplier
    generic map(
            re_multiplicator=>16134, --- 0.984741210938 + j-0.173950195312
            im_multiplicator=>-2850
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1825),
            data_im_in=>first_stage_im_out(1825),
            product_re_out=>mul_re_out(1825),
            product_im_out=>mul_im_out(1825)
        );

    UMUL_1826 : complex_multiplier
    generic map(
            re_multiplicator=>15392, --- 0.939453125 + j-0.342651367188
            im_multiplicator=>-5614
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1826),
            data_im_in=>first_stage_im_out(1826),
            product_re_out=>mul_re_out(1826),
            product_im_out=>mul_im_out(1826)
        );

    UMUL_1827 : complex_multiplier
    generic map(
            re_multiplicator=>14180, --- 0.865478515625 + j-0.500854492188
            im_multiplicator=>-8206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1827),
            data_im_in=>first_stage_im_out(1827),
            product_re_out=>mul_re_out(1827),
            product_im_out=>mul_im_out(1827)
        );

    UMUL_1828 : complex_multiplier
    generic map(
            re_multiplicator=>12536, --- 0.76513671875 + j-0.643798828125
            im_multiplicator=>-10548
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1828),
            data_im_in=>first_stage_im_out(1828),
            product_re_out=>mul_re_out(1828),
            product_im_out=>mul_im_out(1828)
        );

    UMUL_1829 : complex_multiplier
    generic map(
            re_multiplicator=>10510, --- 0.641479492188 + j-0.76708984375
            im_multiplicator=>-12568
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1829),
            data_im_in=>first_stage_im_out(1829),
            product_re_out=>mul_re_out(1829),
            product_im_out=>mul_im_out(1829)
        );

    UMUL_1830 : complex_multiplier
    generic map(
            re_multiplicator=>8162, --- 0.498168945312 + j-0.867004394531
            im_multiplicator=>-14205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1830),
            data_im_in=>first_stage_im_out(1830),
            product_re_out=>mul_re_out(1830),
            product_im_out=>mul_im_out(1830)
        );

    UMUL_1831 : complex_multiplier
    generic map(
            re_multiplicator=>5566, --- 0.339721679688 + j-0.940490722656
            im_multiplicator=>-15409
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1831),
            data_im_in=>first_stage_im_out(1831),
            product_re_out=>mul_re_out(1831),
            product_im_out=>mul_im_out(1831)
        );

    UMUL_1832 : complex_multiplier
    generic map(
            re_multiplicator=>2801, --- 0.170959472656 + j-0.985229492188
            im_multiplicator=>-16142
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1832),
            data_im_in=>first_stage_im_out(1832),
            product_re_out=>mul_re_out(1832),
            product_im_out=>mul_im_out(1832)
        );

    UMUL_1833 : complex_multiplier
    generic map(
            re_multiplicator=>-50, --- -0.0030517578125 + j-0.999938964844
            im_multiplicator=>-16383
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1833),
            data_im_in=>first_stage_im_out(1833),
            product_re_out=>mul_re_out(1833),
            product_im_out=>mul_im_out(1833)
        );

    UMUL_1834 : complex_multiplier
    generic map(
            re_multiplicator=>-2900, --- -0.177001953125 + j-0.984191894531
            im_multiplicator=>-16125
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1834),
            data_im_in=>first_stage_im_out(1834),
            product_re_out=>mul_re_out(1834),
            product_im_out=>mul_im_out(1834)
        );

    UMUL_1835 : complex_multiplier
    generic map(
            re_multiplicator=>-5661, --- -0.345520019531 + j-0.938354492188
            im_multiplicator=>-15374
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1835),
            data_im_in=>first_stage_im_out(1835),
            product_re_out=>mul_re_out(1835),
            product_im_out=>mul_im_out(1835)
        );

    UMUL_1836 : complex_multiplier
    generic map(
            re_multiplicator=>-8249, --- -0.503479003906 + j-0.863952636719
            im_multiplicator=>-14155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1836),
            data_im_in=>first_stage_im_out(1836),
            product_re_out=>mul_re_out(1836),
            product_im_out=>mul_im_out(1836)
        );

    UMUL_1837 : complex_multiplier
    generic map(
            re_multiplicator=>-10586, --- -0.646118164062 + j-0.76318359375
            im_multiplicator=>-12504
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1837),
            data_im_in=>first_stage_im_out(1837),
            product_re_out=>mul_re_out(1837),
            product_im_out=>mul_im_out(1837)
        );

    UMUL_1838 : complex_multiplier
    generic map(
            re_multiplicator=>-12600, --- -0.76904296875 + j-0.639099121094
            im_multiplicator=>-10471
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1838),
            data_im_in=>first_stage_im_out(1838),
            product_re_out=>mul_re_out(1838),
            product_im_out=>mul_im_out(1838)
        );

    UMUL_1839 : complex_multiplier
    generic map(
            re_multiplicator=>-14230, --- -0.868530273438 + j-0.495544433594
            im_multiplicator=>-8119
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1839),
            data_im_in=>first_stage_im_out(1839),
            product_re_out=>mul_re_out(1839),
            product_im_out=>mul_im_out(1839)
        );

    UMUL_1840 : complex_multiplier
    generic map(
            re_multiplicator=>-15426, --- -0.941528320312 + j-0.336853027344
            im_multiplicator=>-5519
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1840),
            data_im_in=>first_stage_im_out(1840),
            product_re_out=>mul_re_out(1840),
            product_im_out=>mul_im_out(1840)
        );

    UMUL_1841 : complex_multiplier
    generic map(
            re_multiplicator=>-16151, --- -0.985778808594 + j-0.167907714844
            im_multiplicator=>-2751
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1841),
            data_im_in=>first_stage_im_out(1841),
            product_re_out=>mul_re_out(1841),
            product_im_out=>mul_im_out(1841)
        );

    UMUL_1842 : complex_multiplier
    generic map(
            re_multiplicator=>-16383, --- -0.999938964844 + j0.006103515625
            im_multiplicator=>100
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1842),
            data_im_in=>first_stage_im_out(1842),
            product_re_out=>mul_re_out(1842),
            product_im_out=>mul_im_out(1842)
        );

    UMUL_1843 : complex_multiplier
    generic map(
            re_multiplicator=>-16116, --- -0.983642578125 + j0.179992675781
            im_multiplicator=>2949
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1843),
            data_im_in=>first_stage_im_out(1843),
            product_re_out=>mul_re_out(1843),
            product_im_out=>mul_im_out(1843)
        );

    UMUL_1844 : complex_multiplier
    generic map(
            re_multiplicator=>-15357, --- -0.937316894531 + j0.348388671875
            im_multiplicator=>5708
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1844),
            data_im_in=>first_stage_im_out(1844),
            product_re_out=>mul_re_out(1844),
            product_im_out=>mul_im_out(1844)
        );

    UMUL_1845 : complex_multiplier
    generic map(
            re_multiplicator=>-14129, --- -0.862365722656 + j0.506164550781
            im_multiplicator=>8293
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1845),
            data_im_in=>first_stage_im_out(1845),
            product_re_out=>mul_re_out(1845),
            product_im_out=>mul_im_out(1845)
        );

    UMUL_1846 : complex_multiplier
    generic map(
            re_multiplicator=>-12471, --- -0.761169433594 + j0.648498535156
            im_multiplicator=>10625
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1846),
            data_im_in=>first_stage_im_out(1846),
            product_re_out=>mul_re_out(1846),
            product_im_out=>mul_im_out(1846)
        );

    UMUL_1847 : complex_multiplier
    generic map(
            re_multiplicator=>-10432, --- -0.63671875 + j0.771057128906
            im_multiplicator=>12633
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1847),
            data_im_in=>first_stage_im_out(1847),
            product_re_out=>mul_re_out(1847),
            product_im_out=>mul_im_out(1847)
        );

    UMUL_1848 : complex_multiplier
    generic map(
            re_multiplicator=>-8075, --- -0.492858886719 + j0.870056152344
            im_multiplicator=>14255
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1848),
            data_im_in=>first_stage_im_out(1848),
            product_re_out=>mul_re_out(1848),
            product_im_out=>mul_im_out(1848)
        );

    UMUL_1849 : complex_multiplier
    generic map(
            re_multiplicator=>-5472, --- -0.333984375 + j0.942565917969
            im_multiplicator=>15443
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1849),
            data_im_in=>first_stage_im_out(1849),
            product_re_out=>mul_re_out(1849),
            product_im_out=>mul_im_out(1849)
        );

    UMUL_1850 : complex_multiplier
    generic map(
            re_multiplicator=>-2701, --- -0.164855957031 + j0.986267089844
            im_multiplicator=>16159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1850),
            data_im_in=>first_stage_im_out(1850),
            product_re_out=>mul_re_out(1850),
            product_im_out=>mul_im_out(1850)
        );

    UMUL_1851 : complex_multiplier
    generic map(
            re_multiplicator=>150, --- 0.0091552734375 + j0.999938964844
            im_multiplicator=>16383
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1851),
            data_im_in=>first_stage_im_out(1851),
            product_re_out=>mul_re_out(1851),
            product_im_out=>mul_im_out(1851)
        );

    UMUL_1852 : complex_multiplier
    generic map(
            re_multiplicator=>2998, --- 0.182983398438 + j0.983093261719
            im_multiplicator=>16107
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1852),
            data_im_in=>first_stage_im_out(1852),
            product_re_out=>mul_re_out(1852),
            product_im_out=>mul_im_out(1852)
        );

    UMUL_1853 : complex_multiplier
    generic map(
            re_multiplicator=>5755, --- 0.351257324219 + j0.936218261719
            im_multiplicator=>15339
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1853),
            data_im_in=>first_stage_im_out(1853),
            product_re_out=>mul_re_out(1853),
            product_im_out=>mul_im_out(1853)
        );

    UMUL_1854 : complex_multiplier
    generic map(
            re_multiplicator=>8336, --- 0.5087890625 + j0.86083984375
            im_multiplicator=>14104
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1854),
            data_im_in=>first_stage_im_out(1854),
            product_re_out=>mul_re_out(1854),
            product_im_out=>mul_im_out(1854)
        );

    UMUL_1855 : complex_multiplier
    generic map(
            re_multiplicator=>10663, --- 0.650817871094 + j0.759155273438
            im_multiplicator=>12438
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1855),
            data_im_in=>first_stage_im_out(1855),
            product_re_out=>mul_re_out(1855),
            product_im_out=>mul_im_out(1855)
        );

    UDELAY_1856_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1856),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1856)
        );
    UDELAY_1856_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1856),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1856)
        );
    USHIFTER_1856_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1856),
            data_out=>mul_re_out(1856)
        );
    USHIFTER_1856_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1856),
            data_out=>mul_im_out(1856)
        );

    UMUL_1857 : complex_multiplier
    generic map(
            re_multiplicator=>16125, --- 0.984191894531 + j-0.177001953125
            im_multiplicator=>-2900
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1857),
            data_im_in=>first_stage_im_out(1857),
            product_re_out=>mul_re_out(1857),
            product_im_out=>mul_im_out(1857)
        );

    UMUL_1858 : complex_multiplier
    generic map(
            re_multiplicator=>15357, --- 0.937316894531 + j-0.348388671875
            im_multiplicator=>-5708
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1858),
            data_im_in=>first_stage_im_out(1858),
            product_re_out=>mul_re_out(1858),
            product_im_out=>mul_im_out(1858)
        );

    UMUL_1859 : complex_multiplier
    generic map(
            re_multiplicator=>14104, --- 0.86083984375 + j-0.5087890625
            im_multiplicator=>-8336
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1859),
            data_im_in=>first_stage_im_out(1859),
            product_re_out=>mul_re_out(1859),
            product_im_out=>mul_im_out(1859)
        );

    UMUL_1860 : complex_multiplier
    generic map(
            re_multiplicator=>12406, --- 0.757202148438 + j-0.653137207031
            im_multiplicator=>-10701
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1860),
            data_im_in=>first_stage_im_out(1860),
            product_re_out=>mul_re_out(1860),
            product_im_out=>mul_im_out(1860)
        );

    UMUL_1861 : complex_multiplier
    generic map(
            re_multiplicator=>10315, --- 0.629577636719 + j-0.77685546875
            im_multiplicator=>-12728
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1861),
            data_im_in=>first_stage_im_out(1861),
            product_re_out=>mul_re_out(1861),
            product_im_out=>mul_im_out(1861)
        );

    UMUL_1862 : complex_multiplier
    generic map(
            re_multiplicator=>7900, --- 0.482177734375 + j-0.876037597656
            im_multiplicator=>-14353
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1862),
            data_im_in=>first_stage_im_out(1862),
            product_re_out=>mul_re_out(1862),
            product_im_out=>mul_im_out(1862)
        );

    UMUL_1863 : complex_multiplier
    generic map(
            re_multiplicator=>5234, --- 0.319458007812 + j-0.947570800781
            im_multiplicator=>-15525
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1863),
            data_im_in=>first_stage_im_out(1863),
            product_re_out=>mul_re_out(1863),
            product_im_out=>mul_im_out(1863)
        );

    UMUL_1864 : complex_multiplier
    generic map(
            re_multiplicator=>2404, --- 0.146728515625 + j-0.989135742188
            im_multiplicator=>-16206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1864),
            data_im_in=>first_stage_im_out(1864),
            product_re_out=>mul_re_out(1864),
            product_im_out=>mul_im_out(1864)
        );

    UMUL_1865 : complex_multiplier
    generic map(
            re_multiplicator=>-502, --- -0.0306396484375 + j-0.99951171875
            im_multiplicator=>-16376
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1865),
            data_im_in=>first_stage_im_out(1865),
            product_re_out=>mul_re_out(1865),
            product_im_out=>mul_im_out(1865)
        );

    UMUL_1866 : complex_multiplier
    generic map(
            re_multiplicator=>-3393, --- -0.207092285156 + j-0.978271484375
            im_multiplicator=>-16028
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1866),
            data_im_in=>first_stage_im_out(1866),
            product_re_out=>mul_re_out(1866),
            product_im_out=>mul_im_out(1866)
        );

    UMUL_1867 : complex_multiplier
    generic map(
            re_multiplicator=>-6176, --- -0.376953125 + j-0.926208496094
            im_multiplicator=>-15175
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1867),
            data_im_in=>first_stage_im_out(1867),
            product_re_out=>mul_re_out(1867),
            product_im_out=>mul_im_out(1867)
        );

    UMUL_1868 : complex_multiplier
    generic map(
            re_multiplicator=>-8765, --- -0.534973144531 + j-0.844848632812
            im_multiplicator=>-13842
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1868),
            data_im_in=>first_stage_im_out(1868),
            product_re_out=>mul_re_out(1868),
            product_im_out=>mul_im_out(1868)
        );

    UMUL_1869 : complex_multiplier
    generic map(
            re_multiplicator=>-11077, --- -0.676086425781 + j-0.73681640625
            im_multiplicator=>-12072
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1869),
            data_im_in=>first_stage_im_out(1869),
            product_re_out=>mul_re_out(1869),
            product_im_out=>mul_im_out(1869)
        );

    UMUL_1870 : complex_multiplier
    generic map(
            re_multiplicator=>-13038, --- -0.795776367188 + j-0.60546875
            im_multiplicator=>-9920
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1870),
            data_im_in=>first_stage_im_out(1870),
            product_re_out=>mul_re_out(1870),
            product_im_out=>mul_im_out(1870)
        );

    UMUL_1871 : complex_multiplier
    generic map(
            re_multiplicator=>-14589, --- -0.890441894531 + j-0.455078125
            im_multiplicator=>-7456
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1871),
            data_im_in=>first_stage_im_out(1871),
            product_re_out=>mul_re_out(1871),
            product_im_out=>mul_im_out(1871)
        );

    UMUL_1872 : complex_multiplier
    generic map(
            re_multiplicator=>-15678, --- -0.956909179688 + j-0.290283203125
            im_multiplicator=>-4756
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1872),
            data_im_in=>first_stage_im_out(1872),
            product_re_out=>mul_re_out(1872),
            product_im_out=>mul_im_out(1872)
        );

    UMUL_1873 : complex_multiplier
    generic map(
            re_multiplicator=>-16272, --- -0.9931640625 + j-0.116271972656
            im_multiplicator=>-1905
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1873),
            data_im_in=>first_stage_im_out(1873),
            product_re_out=>mul_re_out(1873),
            product_im_out=>mul_im_out(1873)
        );

    UMUL_1874 : complex_multiplier
    generic map(
            re_multiplicator=>-16353, --- -0.998107910156 + j0.061279296875
            im_multiplicator=>1004
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1874),
            data_im_in=>first_stage_im_out(1874),
            product_re_out=>mul_re_out(1874),
            product_im_out=>mul_im_out(1874)
        );

    UMUL_1875 : complex_multiplier
    generic map(
            re_multiplicator=>-15917, --- -0.971496582031 + j0.236999511719
            im_multiplicator=>3883
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1875),
            data_im_in=>first_stage_im_out(1875),
            product_re_out=>mul_re_out(1875),
            product_im_out=>mul_im_out(1875)
        );

    UMUL_1876 : complex_multiplier
    generic map(
            re_multiplicator=>-14978, --- -0.914184570312 + j0.405212402344
            im_multiplicator=>6639
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1876),
            data_im_in=>first_stage_im_out(1876),
            product_re_out=>mul_re_out(1876),
            product_im_out=>mul_im_out(1876)
        );

    UMUL_1877 : complex_multiplier
    generic map(
            re_multiplicator=>-13566, --- -0.828002929688 + j0.560607910156
            im_multiplicator=>9185
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1877),
            data_im_in=>first_stage_im_out(1877),
            product_re_out=>mul_re_out(1877),
            product_im_out=>mul_im_out(1877)
        );

    UMUL_1878 : complex_multiplier
    generic map(
            re_multiplicator=>-11726, --- -0.715698242188 + j0.698364257812
            im_multiplicator=>11442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1878),
            data_im_in=>first_stage_im_out(1878),
            product_re_out=>mul_re_out(1878),
            product_im_out=>mul_im_out(1878)
        );

    UMUL_1879 : complex_multiplier
    generic map(
            re_multiplicator=>-9516, --- -0.580810546875 + j0.814025878906
            im_multiplicator=>13337
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1879),
            data_im_in=>first_stage_im_out(1879),
            product_re_out=>mul_re_out(1879),
            product_im_out=>mul_im_out(1879)
        );

    UMUL_1880 : complex_multiplier
    generic map(
            re_multiplicator=>-7005, --- -0.427551269531 + j0.903930664062
            im_multiplicator=>14810
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1880),
            data_im_in=>first_stage_im_out(1880),
            product_re_out=>mul_re_out(1880),
            product_im_out=>mul_im_out(1880)
        );

    UMUL_1881 : complex_multiplier
    generic map(
            re_multiplicator=>-4272, --- -0.2607421875 + j0.965393066406
            im_multiplicator=>15817
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1881),
            data_im_in=>first_stage_im_out(1881),
            product_re_out=>mul_re_out(1881),
            product_im_out=>mul_im_out(1881)
        );

    UMUL_1882 : complex_multiplier
    generic map(
            re_multiplicator=>-1405, --- -0.0857543945312 + j0.996276855469
            im_multiplicator=>16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1882),
            data_im_in=>first_stage_im_out(1882),
            product_re_out=>mul_re_out(1882),
            product_im_out=>mul_im_out(1882)
        );

    UMUL_1883 : complex_multiplier
    generic map(
            re_multiplicator=>1505, --- 0.0918579101562 + j0.995727539062
            im_multiplicator=>16314
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1883),
            data_im_in=>first_stage_im_out(1883),
            product_re_out=>mul_re_out(1883),
            product_im_out=>mul_im_out(1883)
        );

    UMUL_1884 : complex_multiplier
    generic map(
            re_multiplicator=>4369, --- 0.266662597656 + j0.963745117188
            im_multiplicator=>15790
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1884),
            data_im_in=>first_stage_im_out(1884),
            product_re_out=>mul_re_out(1884),
            product_im_out=>mul_im_out(1884)
        );

    UMUL_1885 : complex_multiplier
    generic map(
            re_multiplicator=>7095, --- 0.433044433594 + j0.901306152344
            im_multiplicator=>14767
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1885),
            data_im_in=>first_stage_im_out(1885),
            product_re_out=>mul_re_out(1885),
            product_im_out=>mul_im_out(1885)
        );

    UMUL_1886 : complex_multiplier
    generic map(
            re_multiplicator=>9597, --- 0.585754394531 + j0.810424804688
            im_multiplicator=>13278
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1886),
            data_im_in=>first_stage_im_out(1886),
            product_re_out=>mul_re_out(1886),
            product_im_out=>mul_im_out(1886)
        );

    UMUL_1887 : complex_multiplier
    generic map(
            re_multiplicator=>11796, --- 0.719970703125 + j0.693969726562
            im_multiplicator=>11370
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1887),
            data_im_in=>first_stage_im_out(1887),
            product_re_out=>mul_re_out(1887),
            product_im_out=>mul_im_out(1887)
        );

    UDELAY_1888_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1888),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1888)
        );
    UDELAY_1888_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1888),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1888)
        );
    USHIFTER_1888_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1888),
            data_out=>mul_re_out(1888)
        );
    USHIFTER_1888_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1888),
            data_out=>mul_im_out(1888)
        );

    UMUL_1889 : complex_multiplier
    generic map(
            re_multiplicator=>16116, --- 0.983642578125 + j-0.179992675781
            im_multiplicator=>-2949
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1889),
            data_im_in=>first_stage_im_out(1889),
            product_re_out=>mul_re_out(1889),
            product_im_out=>mul_im_out(1889)
        );

    UMUL_1890 : complex_multiplier
    generic map(
            re_multiplicator=>15322, --- 0.935180664062 + j-0.354125976562
            im_multiplicator=>-5802
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1890),
            data_im_in=>first_stage_im_out(1890),
            product_re_out=>mul_re_out(1890),
            product_im_out=>mul_im_out(1890)
        );

    UMUL_1891 : complex_multiplier
    generic map(
            re_multiplicator=>14027, --- 0.856140136719 + j-0.516723632812
            im_multiplicator=>-8466
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1891),
            data_im_in=>first_stage_im_out(1891),
            product_re_out=>mul_re_out(1891),
            product_im_out=>mul_im_out(1891)
        );

    UMUL_1892 : complex_multiplier
    generic map(
            re_multiplicator=>12273, --- 0.749084472656 + j-0.662414550781
            im_multiplicator=>-10853
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1892),
            data_im_in=>first_stage_im_out(1892),
            product_re_out=>mul_re_out(1892),
            product_im_out=>mul_im_out(1892)
        );

    UMUL_1893 : complex_multiplier
    generic map(
            re_multiplicator=>10119, --- 0.617614746094 + j-0.786437988281
            im_multiplicator=>-12885
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1893),
            data_im_in=>first_stage_im_out(1893),
            product_re_out=>mul_re_out(1893),
            product_im_out=>mul_im_out(1893)
        );

    UMUL_1894 : complex_multiplier
    generic map(
            re_multiplicator=>7634, --- 0.465942382812 + j-0.884765625
            im_multiplicator=>-14496
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1894),
            data_im_in=>first_stage_im_out(1894),
            product_re_out=>mul_re_out(1894),
            product_im_out=>mul_im_out(1894)
        );

    UMUL_1895 : complex_multiplier
    generic map(
            re_multiplicator=>4900, --- 0.299072265625 + j-0.954223632812
            im_multiplicator=>-15634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1895),
            data_im_in=>first_stage_im_out(1895),
            product_re_out=>mul_re_out(1895),
            product_im_out=>mul_im_out(1895)
        );

    UMUL_1896 : complex_multiplier
    generic map(
            re_multiplicator=>2005, --- 0.122375488281 + j-0.992431640625
            im_multiplicator=>-16260
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1896),
            data_im_in=>first_stage_im_out(1896),
            product_re_out=>mul_re_out(1896),
            product_im_out=>mul_im_out(1896)
        );

    UMUL_1897 : complex_multiplier
    generic map(
            re_multiplicator=>-954, --- -0.0582275390625 + j-0.998291015625
            im_multiplicator=>-16356
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1897),
            data_im_in=>first_stage_im_out(1897),
            product_re_out=>mul_re_out(1897),
            product_im_out=>mul_im_out(1897)
        );

    UMUL_1898 : complex_multiplier
    generic map(
            re_multiplicator=>-3883, --- -0.236999511719 + j-0.971496582031
            im_multiplicator=>-15917
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1898),
            data_im_in=>first_stage_im_out(1898),
            product_re_out=>mul_re_out(1898),
            product_im_out=>mul_im_out(1898)
        );

    UMUL_1899 : complex_multiplier
    generic map(
            re_multiplicator=>-6685, --- -0.408020019531 + j-0.912902832031
            im_multiplicator=>-14957
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1899),
            data_im_in=>first_stage_im_out(1899),
            product_re_out=>mul_re_out(1899),
            product_im_out=>mul_im_out(1899)
        );

    UMUL_1900 : complex_multiplier
    generic map(
            re_multiplicator=>-9268, --- -0.565673828125 + j-0.824584960938
            im_multiplicator=>-13510
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1900),
            data_im_in=>first_stage_im_out(1900),
            product_re_out=>mul_re_out(1900),
            product_im_out=>mul_im_out(1900)
        );

    UMUL_1901 : complex_multiplier
    generic map(
            re_multiplicator=>-11549, --- -0.704895019531 + j-0.709228515625
            im_multiplicator=>-11620
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1901),
            data_im_in=>first_stage_im_out(1901),
            product_re_out=>mul_re_out(1901),
            product_im_out=>mul_im_out(1901)
        );

    UMUL_1902 : complex_multiplier
    generic map(
            re_multiplicator=>-13452, --- -0.821044921875 + j-0.570739746094
            im_multiplicator=>-9351
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1902),
            data_im_in=>first_stage_im_out(1902),
            product_re_out=>mul_re_out(1902),
            product_im_out=>mul_im_out(1902)
        );

    UMUL_1903 : complex_multiplier
    generic map(
            re_multiplicator=>-14916, --- -0.910400390625 + j-0.413635253906
            im_multiplicator=>-6777
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1903),
            data_im_in=>first_stage_im_out(1903),
            product_re_out=>mul_re_out(1903),
            product_im_out=>mul_im_out(1903)
        );

    UMUL_1904 : complex_multiplier
    generic map(
            re_multiplicator=>-15892, --- -0.969970703125 + j-0.242919921875
            im_multiplicator=>-3980
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1904),
            data_im_in=>first_stage_im_out(1904),
            product_re_out=>mul_re_out(1904),
            product_im_out=>mul_im_out(1904)
        );

    UMUL_1905 : complex_multiplier
    generic map(
            re_multiplicator=>-16350, --- -0.997924804688 + j-0.0643310546875
            im_multiplicator=>-1054
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1905),
            data_im_in=>first_stage_im_out(1905),
            product_re_out=>mul_re_out(1905),
            product_im_out=>mul_im_out(1905)
        );

    UMUL_1906 : complex_multiplier
    generic map(
            re_multiplicator=>-16272, --- -0.9931640625 + j0.116271972656
            im_multiplicator=>1905
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1906),
            data_im_in=>first_stage_im_out(1906),
            product_re_out=>mul_re_out(1906),
            product_im_out=>mul_im_out(1906)
        );

    UMUL_1907 : complex_multiplier
    generic map(
            re_multiplicator=>-15663, --- -0.955993652344 + j0.293212890625
            im_multiplicator=>4804
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1907),
            data_im_in=>first_stage_im_out(1907),
            product_re_out=>mul_re_out(1907),
            product_im_out=>mul_im_out(1907)
        );

    UMUL_1908 : complex_multiplier
    generic map(
            re_multiplicator=>-14543, --- -0.887634277344 + j0.460510253906
            im_multiplicator=>7545
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1908),
            data_im_in=>first_stage_im_out(1908),
            product_re_out=>mul_re_out(1908),
            product_im_out=>mul_im_out(1908)
        );

    UMUL_1909 : complex_multiplier
    generic map(
            re_multiplicator=>-12947, --- -0.790222167969 + j0.61279296875
            im_multiplicator=>10040
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1909),
            data_im_in=>first_stage_im_out(1909),
            product_re_out=>mul_re_out(1909),
            product_im_out=>mul_im_out(1909)
        );

    UMUL_1910 : complex_multiplier
    generic map(
            re_multiplicator=>-10928, --- -0.6669921875 + j0.745056152344
            im_multiplicator=>12207
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1910),
            data_im_in=>first_stage_im_out(1910),
            product_re_out=>mul_re_out(1910),
            product_im_out=>mul_im_out(1910)
        );

    UMUL_1911 : complex_multiplier
    generic map(
            re_multiplicator=>-8552, --- -0.52197265625 + j0.852905273438
            im_multiplicator=>13974
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1911),
            data_im_in=>first_stage_im_out(1911),
            product_re_out=>mul_re_out(1911),
            product_im_out=>mul_im_out(1911)
        );

    UMUL_1912 : complex_multiplier
    generic map(
            re_multiplicator=>-5896, --- -0.35986328125 + j0.932983398438
            im_multiplicator=>15286
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1912),
            data_im_in=>first_stage_im_out(1912),
            product_re_out=>mul_re_out(1912),
            product_im_out=>mul_im_out(1912)
        );

    UMUL_1913 : complex_multiplier
    generic map(
            re_multiplicator=>-3048, --- -0.18603515625 + j0.982482910156
            im_multiplicator=>16097
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1913),
            data_im_in=>first_stage_im_out(1913),
            product_re_out=>mul_re_out(1913),
            product_im_out=>mul_im_out(1913)
        );

    UMUL_1914 : complex_multiplier
    generic map(
            re_multiplicator=>-100, --- -0.006103515625 + j0.999938964844
            im_multiplicator=>16383
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1914),
            data_im_in=>first_stage_im_out(1914),
            product_re_out=>mul_re_out(1914),
            product_im_out=>mul_im_out(1914)
        );

    UMUL_1915 : complex_multiplier
    generic map(
            re_multiplicator=>2850, --- 0.173950195312 + j0.984741210938
            im_multiplicator=>16134
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1915),
            data_im_in=>first_stage_im_out(1915),
            product_re_out=>mul_re_out(1915),
            product_im_out=>mul_im_out(1915)
        );

    UMUL_1916 : complex_multiplier
    generic map(
            re_multiplicator=>5708, --- 0.348388671875 + j0.937316894531
            im_multiplicator=>15357
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1916),
            data_im_in=>first_stage_im_out(1916),
            product_re_out=>mul_re_out(1916),
            product_im_out=>mul_im_out(1916)
        );

    UMUL_1917 : complex_multiplier
    generic map(
            re_multiplicator=>8379, --- 0.511413574219 + j0.859252929688
            im_multiplicator=>14078
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1917),
            data_im_in=>first_stage_im_out(1917),
            product_re_out=>mul_re_out(1917),
            product_im_out=>mul_im_out(1917)
        );

    UMUL_1918 : complex_multiplier
    generic map(
            re_multiplicator=>10777, --- 0.657775878906 + j0.753173828125
            im_multiplicator=>12340
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1918),
            data_im_in=>first_stage_im_out(1918),
            product_re_out=>mul_re_out(1918),
            product_im_out=>mul_im_out(1918)
        );

    UMUL_1919 : complex_multiplier
    generic map(
            re_multiplicator=>12822, --- 0.782592773438 + j0.622436523438
            im_multiplicator=>10198
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1919),
            data_im_in=>first_stage_im_out(1919),
            product_re_out=>mul_re_out(1919),
            product_im_out=>mul_im_out(1919)
        );

    UDELAY_1920_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1920),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1920)
        );
    UDELAY_1920_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1920),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1920)
        );
    USHIFTER_1920_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1920),
            data_out=>mul_re_out(1920)
        );
    USHIFTER_1920_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1920),
            data_out=>mul_im_out(1920)
        );

    UMUL_1921 : complex_multiplier
    generic map(
            re_multiplicator=>16107, --- 0.983093261719 + j-0.182983398438
            im_multiplicator=>-2998
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1921),
            data_im_in=>first_stage_im_out(1921),
            product_re_out=>mul_re_out(1921),
            product_im_out=>mul_im_out(1921)
        );

    UMUL_1922 : complex_multiplier
    generic map(
            re_multiplicator=>15286, --- 0.932983398438 + j-0.35986328125
            im_multiplicator=>-5896
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1922),
            data_im_in=>first_stage_im_out(1922),
            product_re_out=>mul_re_out(1922),
            product_im_out=>mul_im_out(1922)
        );

    UMUL_1923 : complex_multiplier
    generic map(
            re_multiplicator=>13948, --- 0.851318359375 + j-0.524536132812
            im_multiplicator=>-8594
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1923),
            data_im_in=>first_stage_im_out(1923),
            product_re_out=>mul_re_out(1923),
            product_im_out=>mul_im_out(1923)
        );

    UMUL_1924 : complex_multiplier
    generic map(
            re_multiplicator=>12139, --- 0.740905761719 + j-0.671508789062
            im_multiplicator=>-11002
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1924),
            data_im_in=>first_stage_im_out(1924),
            product_re_out=>mul_re_out(1924),
            product_im_out=>mul_im_out(1924)
        );

    UMUL_1925 : complex_multiplier
    generic map(
            re_multiplicator=>9920, --- 0.60546875 + j-0.795776367188
            im_multiplicator=>-13038
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1925),
            data_im_in=>first_stage_im_out(1925),
            product_re_out=>mul_re_out(1925),
            product_im_out=>mul_im_out(1925)
        );

    UMUL_1926 : complex_multiplier
    generic map(
            re_multiplicator=>7366, --- 0.449584960938 + j-0.893188476562
            im_multiplicator=>-14634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1926),
            data_im_in=>first_stage_im_out(1926),
            product_re_out=>mul_re_out(1926),
            product_im_out=>mul_im_out(1926)
        );

    UMUL_1927 : complex_multiplier
    generic map(
            re_multiplicator=>4563, --- 0.278503417969 + j-0.960388183594
            im_multiplicator=>-15735
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1927),
            data_im_in=>first_stage_im_out(1927),
            product_re_out=>mul_re_out(1927),
            product_im_out=>mul_im_out(1927)
        );

    UMUL_1928 : complex_multiplier
    generic map(
            re_multiplicator=>1605, --- 0.0979614257812 + j-0.995178222656
            im_multiplicator=>-16305
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1928),
            data_im_in=>first_stage_im_out(1928),
            product_re_out=>mul_re_out(1928),
            product_im_out=>mul_im_out(1928)
        );

    UMUL_1929 : complex_multiplier
    generic map(
            re_multiplicator=>-1405, --- -0.0857543945312 + j-0.996276855469
            im_multiplicator=>-16323
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1929),
            data_im_in=>first_stage_im_out(1929),
            product_re_out=>mul_re_out(1929),
            product_im_out=>mul_im_out(1929)
        );

    UMUL_1930 : complex_multiplier
    generic map(
            re_multiplicator=>-4369, --- -0.266662597656 + j-0.963745117188
            im_multiplicator=>-15790
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1930),
            data_im_in=>first_stage_im_out(1930),
            product_re_out=>mul_re_out(1930),
            product_im_out=>mul_im_out(1930)
        );

    UMUL_1931 : complex_multiplier
    generic map(
            re_multiplicator=>-7186, --- -0.438598632812 + j-0.898620605469
            im_multiplicator=>-14723
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1931),
            data_im_in=>first_stage_im_out(1931),
            product_re_out=>mul_re_out(1931),
            product_im_out=>mul_im_out(1931)
        );

    UMUL_1932 : complex_multiplier
    generic map(
            re_multiplicator=>-9759, --- -0.595642089844 + j-0.803161621094
            im_multiplicator=>-13159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1932),
            data_im_in=>first_stage_im_out(1932),
            product_re_out=>mul_re_out(1932),
            product_im_out=>mul_im_out(1932)
        );

    UMUL_1933 : complex_multiplier
    generic map(
            re_multiplicator=>-12003, --- -0.732604980469 + j-0.680541992188
            im_multiplicator=>-11150
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1933),
            data_im_in=>first_stage_im_out(1933),
            product_re_out=>mul_re_out(1933),
            product_im_out=>mul_im_out(1933)
        );

    UMUL_1934 : complex_multiplier
    generic map(
            re_multiplicator=>-13842, --- -0.844848632812 + j-0.534973144531
            im_multiplicator=>-8765
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1934),
            data_im_in=>first_stage_im_out(1934),
            product_re_out=>mul_re_out(1934),
            product_im_out=>mul_im_out(1934)
        );

    UMUL_1935 : complex_multiplier
    generic map(
            re_multiplicator=>-15212, --- -0.928466796875 + j-0.371276855469
            im_multiplicator=>-6083
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1935),
            data_im_in=>first_stage_im_out(1935),
            product_re_out=>mul_re_out(1935),
            product_im_out=>mul_im_out(1935)
        );

    UMUL_1936 : complex_multiplier
    generic map(
            re_multiplicator=>-16069, --- -0.980773925781 + j-0.195068359375
            im_multiplicator=>-3196
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1936),
            data_im_in=>first_stage_im_out(1936),
            product_re_out=>mul_re_out(1936),
            product_im_out=>mul_im_out(1936)
        );

    UMUL_1937 : complex_multiplier
    generic map(
            re_multiplicator=>-16382, --- -0.999877929688 + j-0.0122680664062
            im_multiplicator=>-201
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1937),
            data_im_in=>first_stage_im_out(1937),
            product_re_out=>mul_re_out(1937),
            product_im_out=>mul_im_out(1937)
        );

    UMUL_1938 : complex_multiplier
    generic map(
            re_multiplicator=>-16142, --- -0.985229492188 + j0.170959472656
            im_multiplicator=>2801
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1938),
            data_im_in=>first_stage_im_out(1938),
            product_re_out=>mul_re_out(1938),
            product_im_out=>mul_im_out(1938)
        );

    UMUL_1939 : complex_multiplier
    generic map(
            re_multiplicator=>-15357, --- -0.937316894531 + j0.348388671875
            im_multiplicator=>5708
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1939),
            data_im_in=>first_stage_im_out(1939),
            product_re_out=>mul_re_out(1939),
            product_im_out=>mul_im_out(1939)
        );

    UMUL_1940 : complex_multiplier
    generic map(
            re_multiplicator=>-14053, --- -0.857727050781 + j0.514099121094
            im_multiplicator=>8423
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1940),
            data_im_in=>first_stage_im_out(1940),
            product_re_out=>mul_re_out(1940),
            product_im_out=>mul_im_out(1940)
        );

    UMUL_1941 : complex_multiplier
    generic map(
            re_multiplicator=>-12273, --- -0.749084472656 + j0.662414550781
            im_multiplicator=>10853
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1941),
            data_im_in=>first_stage_im_out(1941),
            product_re_out=>mul_re_out(1941),
            product_im_out=>mul_im_out(1941)
        );

    UMUL_1942 : complex_multiplier
    generic map(
            re_multiplicator=>-10079, --- -0.615173339844 + j0.788330078125
            im_multiplicator=>12916
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1942),
            data_im_in=>first_stage_im_out(1942),
            product_re_out=>mul_re_out(1942),
            product_im_out=>mul_im_out(1942)
        );

    UMUL_1943 : complex_multiplier
    generic map(
            re_multiplicator=>-7545, --- -0.460510253906 + j0.887634277344
            im_multiplicator=>14543
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1943),
            data_im_in=>first_stage_im_out(1943),
            product_re_out=>mul_re_out(1943),
            product_im_out=>mul_im_out(1943)
        );

    UMUL_1944 : complex_multiplier
    generic map(
            re_multiplicator=>-4756, --- -0.290283203125 + j0.956909179688
            im_multiplicator=>15678
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1944),
            data_im_in=>first_stage_im_out(1944),
            product_re_out=>mul_re_out(1944),
            product_im_out=>mul_im_out(1944)
        );

    UMUL_1945 : complex_multiplier
    generic map(
            re_multiplicator=>-1805, --- -0.110168457031 + j0.993896484375
            im_multiplicator=>16284
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1945),
            data_im_in=>first_stage_im_out(1945),
            product_re_out=>mul_re_out(1945),
            product_im_out=>mul_im_out(1945)
        );

    UMUL_1946 : complex_multiplier
    generic map(
            re_multiplicator=>1205, --- 0.0735473632812 + j0.997253417969
            im_multiplicator=>16339
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1946),
            data_im_in=>first_stage_im_out(1946),
            product_re_out=>mul_re_out(1946),
            product_im_out=>mul_im_out(1946)
        );

    UMUL_1947 : complex_multiplier
    generic map(
            re_multiplicator=>4175, --- 0.254821777344 + j0.966918945312
            im_multiplicator=>15842
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1947),
            data_im_in=>first_stage_im_out(1947),
            product_re_out=>mul_re_out(1947),
            product_im_out=>mul_im_out(1947)
        );

    UMUL_1948 : complex_multiplier
    generic map(
            re_multiplicator=>7005, --- 0.427551269531 + j0.903930664062
            im_multiplicator=>14810
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1948),
            data_im_in=>first_stage_im_out(1948),
            product_re_out=>mul_re_out(1948),
            product_im_out=>mul_im_out(1948)
        );

    UMUL_1949 : complex_multiplier
    generic map(
            re_multiplicator=>9597, --- 0.585754394531 + j0.810424804688
            im_multiplicator=>13278
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1949),
            data_im_in=>first_stage_im_out(1949),
            product_re_out=>mul_re_out(1949),
            product_im_out=>mul_im_out(1949)
        );

    UMUL_1950 : complex_multiplier
    generic map(
            re_multiplicator=>11866, --- 0.724243164062 + j0.689514160156
            im_multiplicator=>11297
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1950),
            data_im_in=>first_stage_im_out(1950),
            product_re_out=>mul_re_out(1950),
            product_im_out=>mul_im_out(1950)
        );

    UMUL_1951 : complex_multiplier
    generic map(
            re_multiplicator=>13733, --- 0.838195800781 + j0.545288085938
            im_multiplicator=>8934
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1951),
            data_im_in=>first_stage_im_out(1951),
            product_re_out=>mul_re_out(1951),
            product_im_out=>mul_im_out(1951)
        );

    UDELAY_1952_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1952),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1952)
        );
    UDELAY_1952_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1952),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1952)
        );
    USHIFTER_1952_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1952),
            data_out=>mul_re_out(1952)
        );
    USHIFTER_1952_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1952),
            data_out=>mul_im_out(1952)
        );

    UMUL_1953 : complex_multiplier
    generic map(
            re_multiplicator=>16097, --- 0.982482910156 + j-0.18603515625
            im_multiplicator=>-3048
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1953),
            data_im_in=>first_stage_im_out(1953),
            product_re_out=>mul_re_out(1953),
            product_im_out=>mul_im_out(1953)
        );

    UMUL_1954 : complex_multiplier
    generic map(
            re_multiplicator=>15249, --- 0.930725097656 + j-0.365600585938
            im_multiplicator=>-5990
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1954),
            data_im_in=>first_stage_im_out(1954),
            product_re_out=>mul_re_out(1954),
            product_im_out=>mul_im_out(1954)
        );

    UMUL_1955 : complex_multiplier
    generic map(
            re_multiplicator=>13868, --- 0.846435546875 + j-0.532348632812
            im_multiplicator=>-8722
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1955),
            data_im_in=>first_stage_im_out(1955),
            product_re_out=>mul_re_out(1955),
            product_im_out=>mul_im_out(1955)
        );

    UMUL_1956 : complex_multiplier
    generic map(
            re_multiplicator=>12003, --- 0.732604980469 + j-0.680541992188
            im_multiplicator=>-11150
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1956),
            data_im_in=>first_stage_im_out(1956),
            product_re_out=>mul_re_out(1956),
            product_im_out=>mul_im_out(1956)
        );

    UMUL_1957 : complex_multiplier
    generic map(
            re_multiplicator=>9719, --- 0.593200683594 + j-0.804992675781
            im_multiplicator=>-13189
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1957),
            data_im_in=>first_stage_im_out(1957),
            product_re_out=>mul_re_out(1957),
            product_im_out=>mul_im_out(1957)
        );

    UMUL_1958 : complex_multiplier
    generic map(
            re_multiplicator=>7095, --- 0.433044433594 + j-0.901306152344
            im_multiplicator=>-14767
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1958),
            data_im_in=>first_stage_im_out(1958),
            product_re_out=>mul_re_out(1958),
            product_im_out=>mul_im_out(1958)
        );

    UMUL_1959 : complex_multiplier
    generic map(
            re_multiplicator=>4224, --- 0.2578125 + j-0.966186523438
            im_multiplicator=>-15830
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1959),
            data_im_in=>first_stage_im_out(1959),
            product_re_out=>mul_re_out(1959),
            product_im_out=>mul_im_out(1959)
        );

    UMUL_1960 : complex_multiplier
    generic map(
            re_multiplicator=>1205, --- 0.0735473632812 + j-0.997253417969
            im_multiplicator=>-16339
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1960),
            data_im_in=>first_stage_im_out(1960),
            product_re_out=>mul_re_out(1960),
            product_im_out=>mul_im_out(1960)
        );

    UMUL_1961 : complex_multiplier
    generic map(
            re_multiplicator=>-1855, --- -0.113220214844 + j-0.993530273438
            im_multiplicator=>-16278
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1961),
            data_im_in=>first_stage_im_out(1961),
            product_re_out=>mul_re_out(1961),
            product_im_out=>mul_im_out(1961)
        );

    UMUL_1962 : complex_multiplier
    generic map(
            re_multiplicator=>-4852, --- -0.296142578125 + j-0.955139160156
            im_multiplicator=>-15649
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1962),
            data_im_in=>first_stage_im_out(1962),
            product_re_out=>mul_re_out(1962),
            product_im_out=>mul_im_out(1962)
        );

    UMUL_1963 : complex_multiplier
    generic map(
            re_multiplicator=>-7678, --- -0.468627929688 + j-0.883361816406
            im_multiplicator=>-14473
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1963),
            data_im_in=>first_stage_im_out(1963),
            product_re_out=>mul_re_out(1963),
            product_im_out=>mul_im_out(1963)
        );

    UMUL_1964 : complex_multiplier
    generic map(
            re_multiplicator=>-10237, --- -0.624816894531 + j-0.780700683594
            im_multiplicator=>-12791
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1964),
            data_im_in=>first_stage_im_out(1964),
            product_re_out=>mul_re_out(1964),
            product_im_out=>mul_im_out(1964)
        );

    UMUL_1965 : complex_multiplier
    generic map(
            re_multiplicator=>-12438, --- -0.759155273438 + j-0.650817871094
            im_multiplicator=>-10663
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1965),
            data_im_in=>first_stage_im_out(1965),
            product_re_out=>mul_re_out(1965),
            product_im_out=>mul_im_out(1965)
        );

    UMUL_1966 : complex_multiplier
    generic map(
            re_multiplicator=>-14205, --- -0.867004394531 + j-0.498168945312
            im_multiplicator=>-8162
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1966),
            data_im_in=>first_stage_im_out(1966),
            product_re_out=>mul_re_out(1966),
            product_im_out=>mul_im_out(1966)
        );

    UMUL_1967 : complex_multiplier
    generic map(
            re_multiplicator=>-15476, --- -0.944580078125 + j-0.328186035156
            im_multiplicator=>-5377
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1967),
            data_im_in=>first_stage_im_out(1967),
            product_re_out=>mul_re_out(1967),
            product_im_out=>mul_im_out(1967)
        );

    UMUL_1968 : complex_multiplier
    generic map(
            re_multiplicator=>-16206, --- -0.989135742188 + j-0.146728515625
            im_multiplicator=>-2404
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1968),
            data_im_in=>first_stage_im_out(1968),
            product_re_out=>mul_re_out(1968),
            product_im_out=>mul_im_out(1968)
        );

    UMUL_1969 : complex_multiplier
    generic map(
            re_multiplicator=>-16370, --- -0.999145507812 + j0.0398559570312
            im_multiplicator=>653
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1969),
            data_im_in=>first_stage_im_out(1969),
            product_re_out=>mul_re_out(1969),
            product_im_out=>mul_im_out(1969)
        );

    UMUL_1970 : complex_multiplier
    generic map(
            re_multiplicator=>-15963, --- -0.974304199219 + j0.225036621094
            im_multiplicator=>3687
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1970),
            data_im_in=>first_stage_im_out(1970),
            product_re_out=>mul_re_out(1970),
            product_im_out=>mul_im_out(1970)
        );

    UMUL_1971 : complex_multiplier
    generic map(
            re_multiplicator=>-14998, --- -0.915405273438 + j0.402404785156
            im_multiplicator=>6593
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1971),
            data_im_in=>first_stage_im_out(1971),
            product_re_out=>mul_re_out(1971),
            product_im_out=>mul_im_out(1971)
        );

    UMUL_1972 : complex_multiplier
    generic map(
            re_multiplicator=>-13510, --- -0.824584960938 + j0.565673828125
            im_multiplicator=>9268
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1972),
            data_im_in=>first_stage_im_out(1972),
            product_re_out=>mul_re_out(1972),
            product_im_out=>mul_im_out(1972)
        );

    UMUL_1973 : complex_multiplier
    generic map(
            re_multiplicator=>-11549, --- -0.704895019531 + j0.709228515625
            im_multiplicator=>11620
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1973),
            data_im_in=>first_stage_im_out(1973),
            product_re_out=>mul_re_out(1973),
            product_im_out=>mul_im_out(1973)
        );

    UMUL_1974 : complex_multiplier
    generic map(
            re_multiplicator=>-9185, --- -0.560607910156 + j0.828002929688
            im_multiplicator=>13566
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1974),
            data_im_in=>first_stage_im_out(1974),
            product_re_out=>mul_re_out(1974),
            product_im_out=>mul_im_out(1974)
        );

    UMUL_1975 : complex_multiplier
    generic map(
            re_multiplicator=>-6501, --- -0.396789550781 + j0.917846679688
            im_multiplicator=>15038
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1975),
            data_im_in=>first_stage_im_out(1975),
            product_re_out=>mul_re_out(1975),
            product_im_out=>mul_im_out(1975)
        );

    UMUL_1976 : complex_multiplier
    generic map(
            re_multiplicator=>-3589, --- -0.219055175781 + j0.975646972656
            im_multiplicator=>15985
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1976),
            data_im_in=>first_stage_im_out(1976),
            product_re_out=>mul_re_out(1976),
            product_im_out=>mul_im_out(1976)
        );

    UMUL_1977 : complex_multiplier
    generic map(
            re_multiplicator=>-552, --- -0.03369140625 + j0.999389648438
            im_multiplicator=>16374
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1977),
            data_im_in=>first_stage_im_out(1977),
            product_re_out=>mul_re_out(1977),
            product_im_out=>mul_im_out(1977)
        );

    UMUL_1978 : complex_multiplier
    generic map(
            re_multiplicator=>2503, --- 0.152770996094 + j0.988220214844
            im_multiplicator=>16191
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1978),
            data_im_in=>first_stage_im_out(1978),
            product_re_out=>mul_re_out(1978),
            product_im_out=>mul_im_out(1978)
        );

    UMUL_1979 : complex_multiplier
    generic map(
            re_multiplicator=>5472, --- 0.333984375 + j0.942565917969
            im_multiplicator=>15443
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1979),
            data_im_in=>first_stage_im_out(1979),
            product_re_out=>mul_re_out(1979),
            product_im_out=>mul_im_out(1979)
        );

    UMUL_1980 : complex_multiplier
    generic map(
            re_multiplicator=>8249, --- 0.503479003906 + j0.863952636719
            im_multiplicator=>14155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1980),
            data_im_in=>first_stage_im_out(1980),
            product_re_out=>mul_re_out(1980),
            product_im_out=>mul_im_out(1980)
        );

    UMUL_1981 : complex_multiplier
    generic map(
            re_multiplicator=>10739, --- 0.655456542969 + j0.755187988281
            im_multiplicator=>12373
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1981),
            data_im_in=>first_stage_im_out(1981),
            product_re_out=>mul_re_out(1981),
            product_im_out=>mul_im_out(1981)
        );

    UMUL_1982 : complex_multiplier
    generic map(
            re_multiplicator=>12854, --- 0.784545898438 + j0.620056152344
            im_multiplicator=>10159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1982),
            data_im_in=>first_stage_im_out(1982),
            product_re_out=>mul_re_out(1982),
            product_im_out=>mul_im_out(1982)
        );

    UMUL_1983 : complex_multiplier
    generic map(
            re_multiplicator=>14519, --- 0.886169433594 + j0.463256835938
            im_multiplicator=>7590
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1983),
            data_im_in=>first_stage_im_out(1983),
            product_re_out=>mul_re_out(1983),
            product_im_out=>mul_im_out(1983)
        );

    UDELAY_1984_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(1984),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(1984)
        );
    UDELAY_1984_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(1984),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(1984)
        );
    USHIFTER_1984_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(1984),
            data_out=>mul_re_out(1984)
        );
    USHIFTER_1984_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(1984),
            data_out=>mul_im_out(1984)
        );

    UMUL_1985 : complex_multiplier
    generic map(
            re_multiplicator=>16088, --- 0.98193359375 + j-0.189025878906
            im_multiplicator=>-3097
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1985),
            data_im_in=>first_stage_im_out(1985),
            product_re_out=>mul_re_out(1985),
            product_im_out=>mul_im_out(1985)
        );

    UMUL_1986 : complex_multiplier
    generic map(
            re_multiplicator=>15212, --- 0.928466796875 + j-0.371276855469
            im_multiplicator=>-6083
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1986),
            data_im_in=>first_stage_im_out(1986),
            product_re_out=>mul_re_out(1986),
            product_im_out=>mul_im_out(1986)
        );

    UMUL_1987 : complex_multiplier
    generic map(
            re_multiplicator=>13788, --- 0.841552734375 + j-0.540161132812
            im_multiplicator=>-8850
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1987),
            data_im_in=>first_stage_im_out(1987),
            product_re_out=>mul_re_out(1987),
            product_im_out=>mul_im_out(1987)
        );

    UMUL_1988 : complex_multiplier
    generic map(
            re_multiplicator=>11866, --- 0.724243164062 + j-0.689514160156
            im_multiplicator=>-11297
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1988),
            data_im_in=>first_stage_im_out(1988),
            product_re_out=>mul_re_out(1988),
            product_im_out=>mul_im_out(1988)
        );

    UMUL_1989 : complex_multiplier
    generic map(
            re_multiplicator=>9516, --- 0.580810546875 + j-0.814025878906
            im_multiplicator=>-13337
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1989),
            data_im_in=>first_stage_im_out(1989),
            product_re_out=>mul_re_out(1989),
            product_im_out=>mul_im_out(1989)
        );

    UMUL_1990 : complex_multiplier
    generic map(
            re_multiplicator=>6822, --- 0.416381835938 + j-0.909118652344
            im_multiplicator=>-14895
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1990),
            data_im_in=>first_stage_im_out(1990),
            product_re_out=>mul_re_out(1990),
            product_im_out=>mul_im_out(1990)
        );

    UMUL_1991 : complex_multiplier
    generic map(
            re_multiplicator=>3883, --- 0.236999511719 + j-0.971496582031
            im_multiplicator=>-15917
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1991),
            data_im_in=>first_stage_im_out(1991),
            product_re_out=>mul_re_out(1991),
            product_im_out=>mul_im_out(1991)
        );

    UMUL_1992 : complex_multiplier
    generic map(
            re_multiplicator=>803, --- 0.0490112304688 + j-0.998779296875
            im_multiplicator=>-16364
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1992),
            data_im_in=>first_stage_im_out(1992),
            product_re_out=>mul_re_out(1992),
            product_im_out=>mul_im_out(1992)
        );

    UMUL_1993 : complex_multiplier
    generic map(
            re_multiplicator=>-2304, --- -0.140625 + j-0.990051269531
            im_multiplicator=>-16221
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1993),
            data_im_in=>first_stage_im_out(1993),
            product_re_out=>mul_re_out(1993),
            product_im_out=>mul_im_out(1993)
        );

    UMUL_1994 : complex_multiplier
    generic map(
            re_multiplicator=>-5329, --- -0.325256347656 + j-0.945556640625
            im_multiplicator=>-15492
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1994),
            data_im_in=>first_stage_im_out(1994),
            product_re_out=>mul_re_out(1994),
            product_im_out=>mul_im_out(1994)
        );

    UMUL_1995 : complex_multiplier
    generic map(
            re_multiplicator=>-8162, --- -0.498168945312 + j-0.867004394531
            im_multiplicator=>-14205
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1995),
            data_im_in=>first_stage_im_out(1995),
            product_re_out=>mul_re_out(1995),
            product_im_out=>mul_im_out(1995)
        );

    UMUL_1996 : complex_multiplier
    generic map(
            re_multiplicator=>-10701, --- -0.653137207031 + j-0.757202148438
            im_multiplicator=>-12406
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1996),
            data_im_in=>first_stage_im_out(1996),
            product_re_out=>mul_re_out(1996),
            product_im_out=>mul_im_out(1996)
        );

    UMUL_1997 : complex_multiplier
    generic map(
            re_multiplicator=>-12854, --- -0.784545898438 + j-0.620056152344
            im_multiplicator=>-10159
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1997),
            data_im_in=>first_stage_im_out(1997),
            product_re_out=>mul_re_out(1997),
            product_im_out=>mul_im_out(1997)
        );

    UMUL_1998 : complex_multiplier
    generic map(
            re_multiplicator=>-14543, --- -0.887634277344 + j-0.460510253906
            im_multiplicator=>-7545
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1998),
            data_im_in=>first_stage_im_out(1998),
            product_re_out=>mul_re_out(1998),
            product_im_out=>mul_im_out(1998)
        );

    UMUL_1999 : complex_multiplier
    generic map(
            re_multiplicator=>-15707, --- -0.958679199219 + j-0.284362792969
            im_multiplicator=>-4659
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(1999),
            data_im_in=>first_stage_im_out(1999),
            product_re_out=>mul_re_out(1999),
            product_im_out=>mul_im_out(1999)
        );

    UMUL_2000 : complex_multiplier
    generic map(
            re_multiplicator=>-16305, --- -0.995178222656 + j-0.0979614257812
            im_multiplicator=>-1605
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2000),
            data_im_in=>first_stage_im_out(2000),
            product_re_out=>mul_re_out(2000),
            product_im_out=>mul_im_out(2000)
        );

    UMUL_2001 : complex_multiplier
    generic map(
            re_multiplicator=>-16314, --- -0.995727539062 + j0.0918579101562
            im_multiplicator=>1505
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2001),
            data_im_in=>first_stage_im_out(2001),
            product_re_out=>mul_re_out(2001),
            product_im_out=>mul_im_out(2001)
        );

    UMUL_2002 : complex_multiplier
    generic map(
            re_multiplicator=>-15735, --- -0.960388183594 + j0.278503417969
            im_multiplicator=>4563
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2002),
            data_im_in=>first_stage_im_out(2002),
            product_re_out=>mul_re_out(2002),
            product_im_out=>mul_im_out(2002)
        );

    UMUL_2003 : complex_multiplier
    generic map(
            re_multiplicator=>-14589, --- -0.890441894531 + j0.455078125
            im_multiplicator=>7456
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2003),
            data_im_in=>first_stage_im_out(2003),
            product_re_out=>mul_re_out(2003),
            product_im_out=>mul_im_out(2003)
        );

    UMUL_2004 : complex_multiplier
    generic map(
            re_multiplicator=>-12916, --- -0.788330078125 + j0.615173339844
            im_multiplicator=>10079
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2004),
            data_im_in=>first_stage_im_out(2004),
            product_re_out=>mul_re_out(2004),
            product_im_out=>mul_im_out(2004)
        );

    UMUL_2005 : complex_multiplier
    generic map(
            re_multiplicator=>-10777, --- -0.657775878906 + j0.753173828125
            im_multiplicator=>12340
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2005),
            data_im_in=>first_stage_im_out(2005),
            product_re_out=>mul_re_out(2005),
            product_im_out=>mul_im_out(2005)
        );

    UMUL_2006 : complex_multiplier
    generic map(
            re_multiplicator=>-8249, --- -0.503479003906 + j0.863952636719
            im_multiplicator=>14155
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2006),
            data_im_in=>first_stage_im_out(2006),
            product_re_out=>mul_re_out(2006),
            product_im_out=>mul_im_out(2006)
        );

    UMUL_2007 : complex_multiplier
    generic map(
            re_multiplicator=>-5424, --- -0.3310546875 + j0.943542480469
            im_multiplicator=>15459
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2007),
            data_im_in=>first_stage_im_out(2007),
            product_re_out=>mul_re_out(2007),
            product_im_out=>mul_im_out(2007)
        );

    UMUL_2008 : complex_multiplier
    generic map(
            re_multiplicator=>-2404, --- -0.146728515625 + j0.989135742188
            im_multiplicator=>16206
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2008),
            data_im_in=>first_stage_im_out(2008),
            product_re_out=>mul_re_out(2008),
            product_im_out=>mul_im_out(2008)
        );

    UMUL_2009 : complex_multiplier
    generic map(
            re_multiplicator=>703, --- 0.0429077148438 + j0.9990234375
            im_multiplicator=>16368
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2009),
            data_im_in=>first_stage_im_out(2009),
            product_re_out=>mul_re_out(2009),
            product_im_out=>mul_im_out(2009)
        );

    UMUL_2010 : complex_multiplier
    generic map(
            re_multiplicator=>3785, --- 0.231018066406 + j0.972900390625
            im_multiplicator=>15940
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2010),
            data_im_in=>first_stage_im_out(2010),
            product_re_out=>mul_re_out(2010),
            product_im_out=>mul_im_out(2010)
        );

    UMUL_2011 : complex_multiplier
    generic map(
            re_multiplicator=>6731, --- 0.410827636719 + j0.911682128906
            im_multiplicator=>14937
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2011),
            data_im_in=>first_stage_im_out(2011),
            product_re_out=>mul_re_out(2011),
            product_im_out=>mul_im_out(2011)
        );

    UMUL_2012 : complex_multiplier
    generic map(
            re_multiplicator=>9434, --- 0.575805664062 + j0.817565917969
            im_multiplicator=>13395
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2012),
            data_im_in=>first_stage_im_out(2012),
            product_re_out=>mul_re_out(2012),
            product_im_out=>mul_im_out(2012)
        );

    UMUL_2013 : complex_multiplier
    generic map(
            re_multiplicator=>11796, --- 0.719970703125 + j0.693969726562
            im_multiplicator=>11370
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2013),
            data_im_in=>first_stage_im_out(2013),
            product_re_out=>mul_re_out(2013),
            product_im_out=>mul_im_out(2013)
        );

    UMUL_2014 : complex_multiplier
    generic map(
            re_multiplicator=>13733, --- 0.838195800781 + j0.545288085938
            im_multiplicator=>8934
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2014),
            data_im_in=>first_stage_im_out(2014),
            product_re_out=>mul_re_out(2014),
            product_im_out=>mul_im_out(2014)
        );

    UMUL_2015 : complex_multiplier
    generic map(
            re_multiplicator=>15175, --- 0.926208496094 + j0.376953125
            im_multiplicator=>6176
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2015),
            data_im_in=>first_stage_im_out(2015),
            product_re_out=>mul_re_out(2015),
            product_im_out=>mul_im_out(2015)
        );

    UDELAY_2016_RE : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_re_out(2016),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_re(2016)
        );
    UDELAY_2016_IM : Dff_regN
    generic map(N=>15)
    port map(
            D=>first_stage_im_out(2016),
            clk=>clk,
            ce=>ce,
            rst=>rst,
            Q=>shifter_im(2016)
        );
    USHIFTER_2016_RE: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_re(2016),
            data_out=>mul_re_out(2016)
        );
    USHIFTER_2016_IM: shifter
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_in=>shifter_im(2016),
            data_out=>mul_im_out(2016)
        );

    UMUL_2017 : complex_multiplier
    generic map(
            re_multiplicator=>16078, --- 0.981323242188 + j-0.192077636719
            im_multiplicator=>-3147
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2017),
            data_im_in=>first_stage_im_out(2017),
            product_re_out=>mul_re_out(2017),
            product_im_out=>mul_im_out(2017)
        );

    UMUL_2018 : complex_multiplier
    generic map(
            re_multiplicator=>15175, --- 0.926208496094 + j-0.376953125
            im_multiplicator=>-6176
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2018),
            data_im_in=>first_stage_im_out(2018),
            product_re_out=>mul_re_out(2018),
            product_im_out=>mul_im_out(2018)
        );

    UMUL_2019 : complex_multiplier
    generic map(
            re_multiplicator=>13705, --- 0.836486816406 + j-0.5478515625
            im_multiplicator=>-8976
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2019),
            data_im_in=>first_stage_im_out(2019),
            product_re_out=>mul_re_out(2019),
            product_im_out=>mul_im_out(2019)
        );

    UMUL_2020 : complex_multiplier
    generic map(
            re_multiplicator=>11726, --- 0.715698242188 + j-0.698364257812
            im_multiplicator=>-11442
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2020),
            data_im_in=>first_stage_im_out(2020),
            product_re_out=>mul_re_out(2020),
            product_im_out=>mul_im_out(2020)
        );

    UMUL_2021 : complex_multiplier
    generic map(
            re_multiplicator=>9310, --- 0.568237304688 + j-0.822814941406
            im_multiplicator=>-13481
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2021),
            data_im_in=>first_stage_im_out(2021),
            product_re_out=>mul_re_out(2021),
            product_im_out=>mul_im_out(2021)
        );

    UMUL_2022 : complex_multiplier
    generic map(
            re_multiplicator=>6547, --- 0.399597167969 + j-0.916625976562
            im_multiplicator=>-15018
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2022),
            data_im_in=>first_stage_im_out(2022),
            product_re_out=>mul_re_out(2022),
            product_im_out=>mul_im_out(2022)
        );

    UMUL_2023 : complex_multiplier
    generic map(
            re_multiplicator=>3540, --- 0.216064453125 + j-0.976318359375
            im_multiplicator=>-15996
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2023),
            data_im_in=>first_stage_im_out(2023),
            product_re_out=>mul_re_out(2023),
            product_im_out=>mul_im_out(2023)
        );

    UMUL_2024 : complex_multiplier
    generic map(
            re_multiplicator=>402, --- 0.0245361328125 + j-0.999694824219
            im_multiplicator=>-16379
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2024),
            data_im_in=>first_stage_im_out(2024),
            product_re_out=>mul_re_out(2024),
            product_im_out=>mul_im_out(2024)
        );

    UMUL_2025 : complex_multiplier
    generic map(
            re_multiplicator=>-2751, --- -0.167907714844 + j-0.985778808594
            im_multiplicator=>-16151
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2025),
            data_im_in=>first_stage_im_out(2025),
            product_re_out=>mul_re_out(2025),
            product_im_out=>mul_im_out(2025)
        );

    UMUL_2026 : complex_multiplier
    generic map(
            re_multiplicator=>-5802, --- -0.354125976562 + j-0.935180664062
            im_multiplicator=>-15322
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2026),
            data_im_in=>first_stage_im_out(2026),
            product_re_out=>mul_re_out(2026),
            product_im_out=>mul_im_out(2026)
        );

    UMUL_2027 : complex_multiplier
    generic map(
            re_multiplicator=>-8637, --- -0.527160644531 + j-0.849731445312
            im_multiplicator=>-13922
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2027),
            data_im_in=>first_stage_im_out(2027),
            product_re_out=>mul_re_out(2027),
            product_im_out=>mul_im_out(2027)
        );

    UMUL_2028 : complex_multiplier
    generic map(
            re_multiplicator=>-11150, --- -0.680541992188 + j-0.732604980469
            im_multiplicator=>-12003
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2028),
            data_im_in=>first_stage_im_out(2028),
            product_re_out=>mul_re_out(2028),
            product_im_out=>mul_im_out(2028)
        );

    UMUL_2029 : complex_multiplier
    generic map(
            re_multiplicator=>-13249, --- -0.808654785156 + j-0.588256835938
            im_multiplicator=>-9638
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2029),
            data_im_in=>first_stage_im_out(2029),
            product_re_out=>mul_re_out(2029),
            product_im_out=>mul_im_out(2029)
        );

    UMUL_2030 : complex_multiplier
    generic map(
            re_multiplicator=>-14853, --- -0.906555175781 + j-0.421997070312
            im_multiplicator=>-6914
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2030),
            data_im_in=>first_stage_im_out(2030),
            product_re_out=>mul_re_out(2030),
            product_im_out=>mul_im_out(2030)
        );

    UMUL_2031 : complex_multiplier
    generic map(
            re_multiplicator=>-15905, --- -0.970764160156 + j-0.239990234375
            im_multiplicator=>-3932
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2031),
            data_im_in=>first_stage_im_out(2031),
            product_re_out=>mul_re_out(2031),
            product_im_out=>mul_im_out(2031)
        );

    UMUL_2032 : complex_multiplier
    generic map(
            re_multiplicator=>-16364, --- -0.998779296875 + j-0.0490112304688
            im_multiplicator=>-803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2032),
            data_im_in=>first_stage_im_out(2032),
            product_re_out=>mul_re_out(2032),
            product_im_out=>mul_im_out(2032)
        );

    UMUL_2033 : complex_multiplier
    generic map(
            re_multiplicator=>-16213, --- -0.989562988281 + j0.143676757812
            im_multiplicator=>2354
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2033),
            data_im_in=>first_stage_im_out(2033),
            product_re_out=>mul_re_out(2033),
            product_im_out=>mul_im_out(2033)
        );

    UMUL_2034 : complex_multiplier
    generic map(
            re_multiplicator=>-15459, --- -0.943542480469 + j0.3310546875
            im_multiplicator=>5424
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2034),
            data_im_in=>first_stage_im_out(2034),
            product_re_out=>mul_re_out(2034),
            product_im_out=>mul_im_out(2034)
        );

    UMUL_2035 : complex_multiplier
    generic map(
            re_multiplicator=>-14129, --- -0.862365722656 + j0.506164550781
            im_multiplicator=>8293
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2035),
            data_im_in=>first_stage_im_out(2035),
            product_re_out=>mul_re_out(2035),
            product_im_out=>mul_im_out(2035)
        );

    UMUL_2036 : complex_multiplier
    generic map(
            re_multiplicator=>-12273, --- -0.749084472656 + j0.662414550781
            im_multiplicator=>10853
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2036),
            data_im_in=>first_stage_im_out(2036),
            product_re_out=>mul_re_out(2036),
            product_im_out=>mul_im_out(2036)
        );

    UMUL_2037 : complex_multiplier
    generic map(
            re_multiplicator=>-9960, --- -0.60791015625 + j0.7939453125
            im_multiplicator=>13008
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2037),
            data_im_in=>first_stage_im_out(2037),
            product_re_out=>mul_re_out(2037),
            product_im_out=>mul_im_out(2037)
        );

    UMUL_2038 : complex_multiplier
    generic map(
            re_multiplicator=>-7276, --- -0.444091796875 + j0.895935058594
            im_multiplicator=>14679
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2038),
            data_im_in=>first_stage_im_out(2038),
            product_re_out=>mul_re_out(2038),
            product_im_out=>mul_im_out(2038)
        );

    UMUL_2039 : complex_multiplier
    generic map(
            re_multiplicator=>-4321, --- -0.263732910156 + j0.964538574219
            im_multiplicator=>15803
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2039),
            data_im_in=>first_stage_im_out(2039),
            product_re_out=>mul_re_out(2039),
            product_im_out=>mul_im_out(2039)
        );

    UMUL_2040 : complex_multiplier
    generic map(
            re_multiplicator=>-1205, --- -0.0735473632812 + j0.997253417969
            im_multiplicator=>16339
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2040),
            data_im_in=>first_stage_im_out(2040),
            product_re_out=>mul_re_out(2040),
            product_im_out=>mul_im_out(2040)
        );

    UMUL_2041 : complex_multiplier
    generic map(
            re_multiplicator=>1955, --- 0.119323730469 + j0.992797851562
            im_multiplicator=>16266
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2041),
            data_im_in=>first_stage_im_out(2041),
            product_re_out=>mul_re_out(2041),
            product_im_out=>mul_im_out(2041)
        );

    UMUL_2042 : complex_multiplier
    generic map(
            re_multiplicator=>5043, --- 0.307800292969 + j0.951416015625
            im_multiplicator=>15588
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2042),
            data_im_in=>first_stage_im_out(2042),
            product_re_out=>mul_re_out(2042),
            product_im_out=>mul_im_out(2042)
        );

    UMUL_2043 : complex_multiplier
    generic map(
            re_multiplicator=>7944, --- 0.48486328125 + j0.874572753906
            im_multiplicator=>14329
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2043),
            data_im_in=>first_stage_im_out(2043),
            product_re_out=>mul_re_out(2043),
            product_im_out=>mul_im_out(2043)
        );

    UMUL_2044 : complex_multiplier
    generic map(
            re_multiplicator=>10548, --- 0.643798828125 + j0.76513671875
            im_multiplicator=>12536
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2044),
            data_im_in=>first_stage_im_out(2044),
            product_re_out=>mul_re_out(2044),
            product_im_out=>mul_im_out(2044)
        );

    UMUL_2045 : complex_multiplier
    generic map(
            re_multiplicator=>12760, --- 0.77880859375 + j0.627197265625
            im_multiplicator=>10276
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2045),
            data_im_in=>first_stage_im_out(2045),
            product_re_out=>mul_re_out(2045),
            product_im_out=>mul_im_out(2045)
        );

    UMUL_2046 : complex_multiplier
    generic map(
            re_multiplicator=>14496, --- 0.884765625 + j0.465942382812
            im_multiplicator=>7634
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2046),
            data_im_in=>first_stage_im_out(2046),
            product_re_out=>mul_re_out(2046),
            product_im_out=>mul_im_out(2046)
        );

    UMUL_2047 : complex_multiplier
    generic map(
            re_multiplicator=>15693, --- 0.957824707031 + j0.287292480469
            im_multiplicator=>4707
        )
    port map(
            clk=>clk,
            rst=>rst,
            ce=>ce,
            ctrl=>ctrl_delay,
            data_re_in=>first_stage_re_out(2047),
            data_im_in=>first_stage_im_out(2047),
            product_re_out=>mul_re_out(2047),
            product_im_out=>mul_im_out(2047)
        );

end Behavioral;
